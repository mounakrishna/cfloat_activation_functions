/*
Details:
Has all the common structure, enums used across all the modules in this repo

Author: Mouna Krishna
email: mounakrishna27121999@gmail.com
*/
package types;

  typedef struct {
    Bit#(1) sign; // 1 - Negative, 0 - Positive
    Int#(5) exp;
    Bit#(2) mantissa;
  } cfloat_1_5_2 deriving(Bits, Eq, FShow);

  typedef enum {Tanh, Sigmoid, LeakyReLu, SeLu} Operation deriving(Bits, Eq, FShow);

  typedef struct {
    cfloat_1_5_2 inp;
    Int#(6) bias;
    Operation op;
  } PreprocessStageMeta deriving(Bits, Eq, FShow);

  typedef struct {
    Bit#(1) sign,
    Int#(8) act_exp,
    Bit#(3) act_mantissa,
    Int#(6) bias,
    Operation op;
  } ComputeStageMeta deriving(Bits, Eq, FShow);

  typedef struct {
  } PostprocessStageMeta deriving(Bits, Eq, FShow);

  typedef struct {
    Bit#(1) final_sign,
    Int#(8) final_exp,
    Bit#(3) final_mantissa,
  } OutputStageMeta deriving(Bits, Eq, FShow);

endpackage
