package selu_lut;
  import Vector :: *;
  import FIFOF :: *;
  import GetPut :: *;
  import types :: *;

  interface Ifc_selu_lut_region_1;
    method Tuple2#(Bit#(5), Bit#(2)) mv_sig_output(Bit#(4) exp, Bit#(2) man);
  endinterface

  module mkselu_lut_region_1(Ifc_selu_lut_region_1);
    // range: 42 - 314
    Reg#(Bit#(2)) rg_man_output[220];
    rg_man_output[0] = readOnlyReg(0);
    rg_man_output[1] = readOnlyReg(3);
    rg_man_output[2] = readOnlyReg(3);
    rg_man_output[3] = readOnlyReg(3);
    rg_man_output[4] = readOnlyReg(3);
    rg_man_output[5] = readOnlyReg(3);
    rg_man_output[6] = readOnlyReg(3);
    rg_man_output[7] = readOnlyReg(3);
    rg_man_output[8] = readOnlyReg(3);
    rg_man_output[9] = readOnlyReg(3);
    rg_man_output[10] = readOnlyReg(1);
    rg_man_output[11] = readOnlyReg(1);
    rg_man_output[12] = readOnlyReg(3);
    rg_man_output[13] = readOnlyReg(0);
    rg_man_output[14] = readOnlyReg(1);
    rg_man_output[15] = readOnlyReg(2);
    rg_man_output[16] = readOnlyReg(3);
    rg_man_output[17] = readOnlyReg(0);
    rg_man_output[18] = readOnlyReg(1);
    rg_man_output[19] = readOnlyReg(2);
    rg_man_output[20] = readOnlyReg(3);
    rg_man_output[21] = readOnlyReg(0);
    rg_man_output[22] = readOnlyReg(1);
    rg_man_output[23] = readOnlyReg(2);
    rg_man_output[24] = readOnlyReg(3);
    rg_man_output[25] = readOnlyReg(0);
    rg_man_output[26] = readOnlyReg(1);
    rg_man_output[27] = readOnlyReg(2);
    rg_man_output[28] = readOnlyReg(3);
    rg_man_output[29] = readOnlyReg(0);
    rg_man_output[30] = readOnlyReg(1);
    rg_man_output[31] = readOnlyReg(2);
    rg_man_output[32] = readOnlyReg(3);
    rg_man_output[33] = readOnlyReg(0);
    rg_man_output[34] = readOnlyReg(1);
    rg_man_output[35] = readOnlyReg(2);
    rg_man_output[36] = readOnlyReg(3);
    rg_man_output[37] = readOnlyReg(0);
    rg_man_output[38] = readOnlyReg(1);
    rg_man_output[39] = readOnlyReg(2);
    rg_man_output[40] = readOnlyReg(3);
    rg_man_output[41] = readOnlyReg(0);
    rg_man_output[42] = readOnlyReg(1);
    rg_man_output[43] = readOnlyReg(2);
    rg_man_output[44] = readOnlyReg(3);
    rg_man_output[45] = readOnlyReg(0);
    rg_man_output[46] = readOnlyReg(1);
    rg_man_output[47] = readOnlyReg(2);
    rg_man_output[48] = readOnlyReg(3);
    rg_man_output[49] = readOnlyReg(0);
    rg_man_output[50] = readOnlyReg(1);
    rg_man_output[51] = readOnlyReg(2);
    rg_man_output[52] = readOnlyReg(3);
    rg_man_output[53] = readOnlyReg(0);
    rg_man_output[54] = readOnlyReg(1);
    rg_man_output[55] = readOnlyReg(2);
    rg_man_output[56] = readOnlyReg(3);
    rg_man_output[57] = readOnlyReg(0);
    rg_man_output[58] = readOnlyReg(1);
    rg_man_output[59] = readOnlyReg(2);
    rg_man_output[60] = readOnlyReg(3);
    rg_man_output[61] = readOnlyReg(0);
    rg_man_output[62] = readOnlyReg(1);
    rg_man_output[63] = readOnlyReg(2);
    rg_man_output[64] = readOnlyReg(3);
    rg_man_output[65] = readOnlyReg(0);
    rg_man_output[66] = readOnlyReg(1);
    rg_man_output[67] = readOnlyReg(2);
    rg_man_output[68] = readOnlyReg(3);
    rg_man_output[69] = readOnlyReg(0);
    rg_man_output[70] = readOnlyReg(1);
    rg_man_output[71] = readOnlyReg(2);
    rg_man_output[72] = readOnlyReg(3);
    rg_man_output[73] = readOnlyReg(0);
    rg_man_output[74] = readOnlyReg(1);
    rg_man_output[75] = readOnlyReg(2);
    rg_man_output[76] = readOnlyReg(3);
    rg_man_output[77] = readOnlyReg(0);
    rg_man_output[78] = readOnlyReg(1);
    rg_man_output[79] = readOnlyReg(2);
    rg_man_output[80] = readOnlyReg(3);
    rg_man_output[81] = readOnlyReg(0);
    rg_man_output[82] = readOnlyReg(1);
    rg_man_output[83] = readOnlyReg(2);
    rg_man_output[84] = readOnlyReg(3);
    rg_man_output[85] = readOnlyReg(0);
    rg_man_output[86] = readOnlyReg(1);
    rg_man_output[87] = readOnlyReg(2);
    rg_man_output[88] = readOnlyReg(3);
    rg_man_output[89] = readOnlyReg(0);
    rg_man_output[90] = readOnlyReg(1);
    rg_man_output[91] = readOnlyReg(2);
    rg_man_output[92] = readOnlyReg(3);
    rg_man_output[93] = readOnlyReg(0);
    rg_man_output[94] = readOnlyReg(1);
    rg_man_output[95] = readOnlyReg(2);
    rg_man_output[96] = readOnlyReg(3);
    rg_man_output[97] = readOnlyReg(0);
    rg_man_output[98] = readOnlyReg(1);
    rg_man_output[99] = readOnlyReg(2);
    rg_man_output[100] = readOnlyReg(3);
    rg_man_output[101] = readOnlyReg(0);
    rg_man_output[102] = readOnlyReg(1);
    rg_man_output[103] = readOnlyReg(2);
    rg_man_output[104] = readOnlyReg(3);
    rg_man_output[105] = readOnlyReg(0);
    rg_man_output[106] = readOnlyReg(1);
    rg_man_output[107] = readOnlyReg(2);
    rg_man_output[108] = readOnlyReg(3);
    rg_man_output[109] = readOnlyReg(0);
    rg_man_output[110] = readOnlyReg(1);
    rg_man_output[111] = readOnlyReg(2);
    rg_man_output[112] = readOnlyReg(3);
    rg_man_output[113] = readOnlyReg(0);
    rg_man_output[114] = readOnlyReg(1);
    rg_man_output[115] = readOnlyReg(2);
    rg_man_output[116] = readOnlyReg(3);
    rg_man_output[117] = readOnlyReg(0);
    rg_man_output[118] = readOnlyReg(1);
    rg_man_output[119] = readOnlyReg(2);
    rg_man_output[120] = readOnlyReg(3);
    rg_man_output[121] = readOnlyReg(0);
    rg_man_output[122] = readOnlyReg(1);
    rg_man_output[123] = readOnlyReg(2);
    rg_man_output[124] = readOnlyReg(3);
    rg_man_output[125] = readOnlyReg(0);
    rg_man_output[126] = readOnlyReg(1);
    rg_man_output[127] = readOnlyReg(2);
    rg_man_output[128] = readOnlyReg(3);
    rg_man_output[129] = readOnlyReg(0);
    rg_man_output[130] = readOnlyReg(1);
    rg_man_output[131] = readOnlyReg(2);
    rg_man_output[132] = readOnlyReg(3);
    rg_man_output[133] = readOnlyReg(0);
    rg_man_output[134] = readOnlyReg(1);
    rg_man_output[135] = readOnlyReg(2);
    rg_man_output[136] = readOnlyReg(3);
    rg_man_output[137] = readOnlyReg(0);
    rg_man_output[138] = readOnlyReg(1);
    rg_man_output[139] = readOnlyReg(2);
    rg_man_output[140] = readOnlyReg(3);
    rg_man_output[141] = readOnlyReg(0);
    rg_man_output[142] = readOnlyReg(1);
    rg_man_output[143] = readOnlyReg(2);
    rg_man_output[144] = readOnlyReg(3);
    rg_man_output[145] = readOnlyReg(0);
    rg_man_output[146] = readOnlyReg(1);
    rg_man_output[147] = readOnlyReg(2);
    rg_man_output[148] = readOnlyReg(3);
    rg_man_output[149] = readOnlyReg(0);
    rg_man_output[150] = readOnlyReg(1);
    rg_man_output[151] = readOnlyReg(2);
    rg_man_output[152] = readOnlyReg(3);
    rg_man_output[153] = readOnlyReg(0);
    rg_man_output[154] = readOnlyReg(1);
    rg_man_output[155] = readOnlyReg(2);
    rg_man_output[156] = readOnlyReg(3);
    rg_man_output[157] = readOnlyReg(0);
    rg_man_output[158] = readOnlyReg(1);
    rg_man_output[159] = readOnlyReg(2);
    rg_man_output[160] = readOnlyReg(3);
    rg_man_output[161] = readOnlyReg(0);
    rg_man_output[162] = readOnlyReg(1);
    rg_man_output[163] = readOnlyReg(2);
    rg_man_output[164] = readOnlyReg(3);
    rg_man_output[165] = readOnlyReg(0);
    rg_man_output[166] = readOnlyReg(1);
    rg_man_output[167] = readOnlyReg(2);
    rg_man_output[168] = readOnlyReg(3);
    rg_man_output[169] = readOnlyReg(0);
    rg_man_output[170] = readOnlyReg(1);
    rg_man_output[171] = readOnlyReg(2);
    rg_man_output[172] = readOnlyReg(3);
    rg_man_output[173] = readOnlyReg(0);
    rg_man_output[174] = readOnlyReg(1);
    rg_man_output[175] = readOnlyReg(2);
    rg_man_output[176] = readOnlyReg(3);
    rg_man_output[177] = readOnlyReg(0);
    rg_man_output[178] = readOnlyReg(1);
    rg_man_output[179] = readOnlyReg(2);
    rg_man_output[180] = readOnlyReg(3);
    rg_man_output[181] = readOnlyReg(0);
    rg_man_output[182] = readOnlyReg(1);
    rg_man_output[183] = readOnlyReg(2);
    rg_man_output[184] = readOnlyReg(3);
    rg_man_output[185] = readOnlyReg(0);
    rg_man_output[186] = readOnlyReg(1);
    rg_man_output[187] = readOnlyReg(2);
    rg_man_output[188] = readOnlyReg(3);
    rg_man_output[189] = readOnlyReg(0);
    rg_man_output[190] = readOnlyReg(1);
    rg_man_output[191] = readOnlyReg(2);
    rg_man_output[192] = readOnlyReg(3);
    rg_man_output[193] = readOnlyReg(0);
    rg_man_output[194] = readOnlyReg(1);
    rg_man_output[195] = readOnlyReg(2);
    rg_man_output[196] = readOnlyReg(3);
    rg_man_output[197] = readOnlyReg(0);
    rg_man_output[198] = readOnlyReg(1);
    rg_man_output[199] = readOnlyReg(2);
    rg_man_output[200] = readOnlyReg(3);
    rg_man_output[201] = readOnlyReg(0);
    rg_man_output[202] = readOnlyReg(1);
    rg_man_output[203] = readOnlyReg(2);
    rg_man_output[204] = readOnlyReg(3);
    rg_man_output[205] = readOnlyReg(0);
    rg_man_output[206] = readOnlyReg(1);
    rg_man_output[207] = readOnlyReg(2);
    rg_man_output[208] = readOnlyReg(2);
    rg_man_output[209] = readOnlyReg(0);
    rg_man_output[210] = readOnlyReg(0);
    rg_man_output[211] = readOnlyReg(1);
    rg_man_output[212] = readOnlyReg(2);
    rg_man_output[213] = readOnlyReg(3);
    rg_man_output[214] = readOnlyReg(3);
    rg_man_output[215] = readOnlyReg(3);
    rg_man_output[216] = readOnlyReg(0);
    rg_man_output[217] = readOnlyReg(2);
    rg_man_output[218] = readOnlyReg(2);
    rg_man_output[219] = readOnlyReg(3);
    

    Reg#(Int#(5)) rg_exp_output[220];
    rg_exp_output[0] = readOnlyReg(0);
    rg_exp_output[1] = readOnlyReg(-53);
    rg_exp_output[2] = readOnlyReg(-53);
    rg_exp_output[3] = readOnlyReg(-53);
    rg_exp_output[4] = readOnlyReg(-53);
    rg_exp_output[5] = readOnlyReg(-53);
    rg_exp_output[6] = readOnlyReg(-53);
    rg_exp_output[7] = readOnlyReg(-52);
    rg_exp_output[8] = readOnlyReg(-52);
    rg_exp_output[9] = readOnlyReg(-52);
    rg_exp_output[10] = readOnlyReg(-51);
    rg_exp_output[11] = readOnlyReg(-51);
    rg_exp_output[12] = readOnlyReg(-51);
    rg_exp_output[13] = readOnlyReg(-50);
    rg_exp_output[14] = readOnlyReg(-50);
    rg_exp_output[15] = readOnlyReg(-50);
    rg_exp_output[16] = readOnlyReg(-50);
    rg_exp_output[17] = readOnlyReg(-49);
    rg_exp_output[18] = readOnlyReg(-49);
    rg_exp_output[19] = readOnlyReg(-49);
    rg_exp_output[20] = readOnlyReg(-49);
    rg_exp_output[21] = readOnlyReg(-48);
    rg_exp_output[22] = readOnlyReg(-48);
    rg_exp_output[23] = readOnlyReg(-48);
    rg_exp_output[24] = readOnlyReg(-48);
    rg_exp_output[25] = readOnlyReg(-47);
    rg_exp_output[26] = readOnlyReg(-47);
    rg_exp_output[27] = readOnlyReg(-47);
    rg_exp_output[28] = readOnlyReg(-47);
    rg_exp_output[29] = readOnlyReg(-46);
    rg_exp_output[30] = readOnlyReg(-46);
    rg_exp_output[31] = readOnlyReg(-46);
    rg_exp_output[32] = readOnlyReg(-46);
    rg_exp_output[33] = readOnlyReg(-45);
    rg_exp_output[34] = readOnlyReg(-45);
    rg_exp_output[35] = readOnlyReg(-45);
    rg_exp_output[36] = readOnlyReg(-45);
    rg_exp_output[37] = readOnlyReg(-44);
    rg_exp_output[38] = readOnlyReg(-44);
    rg_exp_output[39] = readOnlyReg(-44);
    rg_exp_output[40] = readOnlyReg(-44);
    rg_exp_output[41] = readOnlyReg(-43);
    rg_exp_output[42] = readOnlyReg(-43);
    rg_exp_output[43] = readOnlyReg(-43);
    rg_exp_output[44] = readOnlyReg(-43);
    rg_exp_output[45] = readOnlyReg(-42);
    rg_exp_output[46] = readOnlyReg(-42);
    rg_exp_output[47] = readOnlyReg(-42);
    rg_exp_output[48] = readOnlyReg(-42);
    rg_exp_output[49] = readOnlyReg(-41);
    rg_exp_output[50] = readOnlyReg(-41);
    rg_exp_output[51] = readOnlyReg(-41);
    rg_exp_output[52] = readOnlyReg(-41);
    rg_exp_output[53] = readOnlyReg(-40);
    rg_exp_output[54] = readOnlyReg(-40);
    rg_exp_output[55] = readOnlyReg(-40);
    rg_exp_output[56] = readOnlyReg(-40);
    rg_exp_output[57] = readOnlyReg(-39);
    rg_exp_output[58] = readOnlyReg(-39);
    rg_exp_output[59] = readOnlyReg(-39);
    rg_exp_output[60] = readOnlyReg(-39);
    rg_exp_output[61] = readOnlyReg(-38);
    rg_exp_output[62] = readOnlyReg(-38);
    rg_exp_output[63] = readOnlyReg(-38);
    rg_exp_output[64] = readOnlyReg(-38);
    rg_exp_output[65] = readOnlyReg(-37);
    rg_exp_output[66] = readOnlyReg(-37);
    rg_exp_output[67] = readOnlyReg(-37);
    rg_exp_output[68] = readOnlyReg(-37);
    rg_exp_output[69] = readOnlyReg(-36);
    rg_exp_output[70] = readOnlyReg(-36);
    rg_exp_output[71] = readOnlyReg(-36);
    rg_exp_output[72] = readOnlyReg(-36);
    rg_exp_output[73] = readOnlyReg(-35);
    rg_exp_output[74] = readOnlyReg(-35);
    rg_exp_output[75] = readOnlyReg(-35);
    rg_exp_output[76] = readOnlyReg(-35);
    rg_exp_output[77] = readOnlyReg(-34);
    rg_exp_output[78] = readOnlyReg(-34);
    rg_exp_output[79] = readOnlyReg(-34);
    rg_exp_output[80] = readOnlyReg(-34);
    rg_exp_output[81] = readOnlyReg(-33);
    rg_exp_output[82] = readOnlyReg(-33);
    rg_exp_output[83] = readOnlyReg(-33);
    rg_exp_output[84] = readOnlyReg(-33);
    rg_exp_output[85] = readOnlyReg(-32);
    rg_exp_output[86] = readOnlyReg(-32);
    rg_exp_output[87] = readOnlyReg(-32);
    rg_exp_output[88] = readOnlyReg(-32);
    rg_exp_output[89] = readOnlyReg(-31);
    rg_exp_output[90] = readOnlyReg(-31);
    rg_exp_output[91] = readOnlyReg(-31);
    rg_exp_output[92] = readOnlyReg(-31);
    rg_exp_output[93] = readOnlyReg(-30);
    rg_exp_output[94] = readOnlyReg(-30);
    rg_exp_output[95] = readOnlyReg(-30);
    rg_exp_output[96] = readOnlyReg(-30);
    rg_exp_output[97] = readOnlyReg(-29);
    rg_exp_output[98] = readOnlyReg(-29);
    rg_exp_output[99] = readOnlyReg(-29);
    rg_exp_output[100] = readOnlyReg(-29);
    rg_exp_output[101] = readOnlyReg(-28);
    rg_exp_output[102] = readOnlyReg(-28);
    rg_exp_output[103] = readOnlyReg(-28);
    rg_exp_output[104] = readOnlyReg(-28);
    rg_exp_output[105] = readOnlyReg(-27);
    rg_exp_output[106] = readOnlyReg(-27);
    rg_exp_output[107] = readOnlyReg(-27);
    rg_exp_output[108] = readOnlyReg(-27);
    rg_exp_output[109] = readOnlyReg(-26);
    rg_exp_output[110] = readOnlyReg(-26);
    rg_exp_output[111] = readOnlyReg(-26);
    rg_exp_output[112] = readOnlyReg(-26);
    rg_exp_output[113] = readOnlyReg(-25);
    rg_exp_output[114] = readOnlyReg(-25);
    rg_exp_output[115] = readOnlyReg(-25);
    rg_exp_output[116] = readOnlyReg(-25);
    rg_exp_output[117] = readOnlyReg(-24);
    rg_exp_output[118] = readOnlyReg(-24);
    rg_exp_output[119] = readOnlyReg(-24);
    rg_exp_output[120] = readOnlyReg(-24);
    rg_exp_output[121] = readOnlyReg(-23);
    rg_exp_output[122] = readOnlyReg(-23);
    rg_exp_output[123] = readOnlyReg(-23);
    rg_exp_output[124] = readOnlyReg(-23);
    rg_exp_output[125] = readOnlyReg(-22);
    rg_exp_output[126] = readOnlyReg(-22);
    rg_exp_output[127] = readOnlyReg(-22);
    rg_exp_output[128] = readOnlyReg(-22);
    rg_exp_output[129] = readOnlyReg(-21);
    rg_exp_output[130] = readOnlyReg(-21);
    rg_exp_output[131] = readOnlyReg(-21);
    rg_exp_output[132] = readOnlyReg(-21);
    rg_exp_output[133] = readOnlyReg(-20);
    rg_exp_output[134] = readOnlyReg(-20);
    rg_exp_output[135] = readOnlyReg(-20);
    rg_exp_output[136] = readOnlyReg(-20);
    rg_exp_output[137] = readOnlyReg(-19);
    rg_exp_output[138] = readOnlyReg(-19);
    rg_exp_output[139] = readOnlyReg(-19);
    rg_exp_output[140] = readOnlyReg(-19);
    rg_exp_output[141] = readOnlyReg(-18);
    rg_exp_output[142] = readOnlyReg(-18);
    rg_exp_output[143] = readOnlyReg(-18);
    rg_exp_output[144] = readOnlyReg(-18);
    rg_exp_output[145] = readOnlyReg(-17);
    rg_exp_output[146] = readOnlyReg(-17);
    rg_exp_output[147] = readOnlyReg(-17);
    rg_exp_output[148] = readOnlyReg(-17);
    rg_exp_output[149] = readOnlyReg(-16);
    rg_exp_output[150] = readOnlyReg(-16);
    rg_exp_output[151] = readOnlyReg(-16);
    rg_exp_output[152] = readOnlyReg(-16);
    rg_exp_output[153] = readOnlyReg(-15);
    rg_exp_output[154] = readOnlyReg(-15);
    rg_exp_output[155] = readOnlyReg(-15);
    rg_exp_output[156] = readOnlyReg(-15);
    rg_exp_output[157] = readOnlyReg(-14);
    rg_exp_output[158] = readOnlyReg(-14);
    rg_exp_output[159] = readOnlyReg(-14);
    rg_exp_output[160] = readOnlyReg(-14);
    rg_exp_output[161] = readOnlyReg(-13);
    rg_exp_output[162] = readOnlyReg(-13);
    rg_exp_output[163] = readOnlyReg(-13);
    rg_exp_output[164] = readOnlyReg(-13);
    rg_exp_output[165] = readOnlyReg(-12);
    rg_exp_output[166] = readOnlyReg(-12);
    rg_exp_output[167] = readOnlyReg(-12);
    rg_exp_output[168] = readOnlyReg(-12);
    rg_exp_output[169] = readOnlyReg(-11);
    rg_exp_output[170] = readOnlyReg(-11);
    rg_exp_output[171] = readOnlyReg(-11);
    rg_exp_output[172] = readOnlyReg(-11);
    rg_exp_output[173] = readOnlyReg(-10);
    rg_exp_output[174] = readOnlyReg(-10);
    rg_exp_output[175] = readOnlyReg(-10);
    rg_exp_output[176] = readOnlyReg(-10);
    rg_exp_output[177] = readOnlyReg(-9);
    rg_exp_output[178] = readOnlyReg(-9);
    rg_exp_output[179] = readOnlyReg(-9);
    rg_exp_output[180] = readOnlyReg(-9);
    rg_exp_output[181] = readOnlyReg(-8);
    rg_exp_output[182] = readOnlyReg(-8);
    rg_exp_output[183] = readOnlyReg(-8);
    rg_exp_output[184] = readOnlyReg(-8);
    rg_exp_output[185] = readOnlyReg(-7);
    rg_exp_output[186] = readOnlyReg(-7);
    rg_exp_output[187] = readOnlyReg(-7);
    rg_exp_output[188] = readOnlyReg(-7);
    rg_exp_output[189] = readOnlyReg(-6);
    rg_exp_output[190] = readOnlyReg(-6);
    rg_exp_output[191] = readOnlyReg(-6);
    rg_exp_output[192] = readOnlyReg(-6);
    rg_exp_output[193] = readOnlyReg(-5);
    rg_exp_output[194] = readOnlyReg(-5);
    rg_exp_output[195] = readOnlyReg(-5);
    rg_exp_output[196] = readOnlyReg(-5);
    rg_exp_output[197] = readOnlyReg(-4);
    rg_exp_output[198] = readOnlyReg(-4);
    rg_exp_output[199] = readOnlyReg(-4);
    rg_exp_output[200] = readOnlyReg(-4);
    rg_exp_output[201] = readOnlyReg(-3);
    rg_exp_output[202] = readOnlyReg(-3);
    rg_exp_output[203] = readOnlyReg(-3);
    rg_exp_output[204] = readOnlyReg(-3);
    rg_exp_output[205] = readOnlyReg(-2);
    rg_exp_output[206] = readOnlyReg(-2);
    rg_exp_output[207] = readOnlyReg(-2);
    rg_exp_output[208] = readOnlyReg(-2);
    rg_exp_output[209] = readOnlyReg(-1);
    rg_exp_output[210] = readOnlyReg(-1);
    rg_exp_output[211] = readOnlyReg(-1);
    rg_exp_output[212] = readOnlyReg(-1);
    rg_exp_output[213] = readOnlyReg(-1);
    rg_exp_output[214] = readOnlyReg(-1);
    rg_exp_output[215] = readOnlyReg(0);
    rg_exp_output[216] = readOnlyReg(0);
    rg_exp_output[217] = readOnlyReg(-2);
    rg_exp_output[218] = readOnlyReg(-1);
    rg_exp_output[219] = readOnlyReg(-1);

    method Tuple2#(Bit#(5), Bit#(2)) mv_sig_output(Bit#(4) exp, Bit#(2) man);
      Bit#(6) index = {man, exp};
      return tuple2(rg_man_output[index], rg_exp_output[index]);
    endmethod
  endmodule

  interface Ifc_selu_lut_region_2;
    method Tuple2#(Bit#(5), Bit#(2)) mv_sig_output(Bit#(4) exp, Bit#(2) man);
  endinterface

  module mkselu_lut_region_2(Ifc_selu_lut_region_2);
    Reg#(Bit#(2)) rg_man_output[376];
    rg_man_output[0] = readOnlyReg(0);
    rg_man_output[1] = readOnlyReg(1);
    rg_man_output[2] = readOnlyReg(2);
    rg_man_output[3] = readOnlyReg(3);
    rg_man_output[4] = readOnlyReg(0);
    rg_man_output[5] = readOnlyReg(1);
    rg_man_output[6] = readOnlyReg(2);
    rg_man_output[7] = readOnlyReg(3);
    rg_man_output[8] = readOnlyReg(0);
    rg_man_output[9] = readOnlyReg(1);
    rg_man_output[10] = readOnlyReg(2);
    rg_man_output[11] = readOnlyReg(3);
    rg_man_output[12] = readOnlyReg(0);
    rg_man_output[13] = readOnlyReg(1);
    rg_man_output[14] = readOnlyReg(2);
    rg_man_output[15] = readOnlyReg(3);
    rg_man_output[16] = readOnlyReg(0);
    rg_man_output[17] = readOnlyReg(1);
    rg_man_output[18] = readOnlyReg(2);
    rg_man_output[19] = readOnlyReg(3);
    rg_man_output[20] = readOnlyReg(0);
    rg_man_output[21] = readOnlyReg(1);
    rg_man_output[22] = readOnlyReg(2);
    rg_man_output[23] = readOnlyReg(3);
    rg_man_output[24] = readOnlyReg(0);
    rg_man_output[25] = readOnlyReg(1);
    rg_man_output[26] = readOnlyReg(2);
    rg_man_output[27] = readOnlyReg(3);
    rg_man_output[28] = readOnlyReg(0);
    rg_man_output[29] = readOnlyReg(1);
    rg_man_output[30] = readOnlyReg(2);
    rg_man_output[31] = readOnlyReg(3);
    rg_man_output[32] = readOnlyReg(0);
    rg_man_output[33] = readOnlyReg(1);
    rg_man_output[34] = readOnlyReg(2);
    rg_man_output[35] = readOnlyReg(3);
    rg_man_output[36] = readOnlyReg(0);
    rg_man_output[37] = readOnlyReg(1);
    rg_man_output[38] = readOnlyReg(2);
    rg_man_output[39] = readOnlyReg(3);
    rg_man_output[40] = readOnlyReg(0);
    rg_man_output[41] = readOnlyReg(1);
    rg_man_output[42] = readOnlyReg(2);
    rg_man_output[43] = readOnlyReg(3);
    rg_man_output[44] = readOnlyReg(0);
    rg_man_output[45] = readOnlyReg(1);
    rg_man_output[46] = readOnlyReg(2);
    rg_man_output[47] = readOnlyReg(3);
    rg_man_output[48] = readOnlyReg(0);
    rg_man_output[49] = readOnlyReg(1);
    rg_man_output[50] = readOnlyReg(2);
    rg_man_output[51] = readOnlyReg(3);
    rg_man_output[52] = readOnlyReg(0);
    rg_man_output[53] = readOnlyReg(1);
    rg_man_output[54] = readOnlyReg(2);
    rg_man_output[55] = readOnlyReg(3);
    rg_man_output[56] = readOnlyReg(0);
    rg_man_output[57] = readOnlyReg(1);
    rg_man_output[58] = readOnlyReg(2);
    rg_man_output[59] = readOnlyReg(3);
    rg_man_output[60] = readOnlyReg(0);
    rg_man_output[61] = readOnlyReg(1);
    rg_man_output[62] = readOnlyReg(2);
    rg_man_output[63] = readOnlyReg(3);
    rg_man_output[64] = readOnlyReg(0);
    rg_man_output[65] = readOnlyReg(1);
    rg_man_output[66] = readOnlyReg(2);
    rg_man_output[67] = readOnlyReg(3);
    rg_man_output[68] = readOnlyReg(0);
    rg_man_output[69] = readOnlyReg(1);
    rg_man_output[70] = readOnlyReg(2);
    rg_man_output[71] = readOnlyReg(3);
    rg_man_output[72] = readOnlyReg(0);
    rg_man_output[73] = readOnlyReg(1);
    rg_man_output[74] = readOnlyReg(2);
    rg_man_output[75] = readOnlyReg(3);
    rg_man_output[76] = readOnlyReg(0);
    rg_man_output[77] = readOnlyReg(1);
    rg_man_output[78] = readOnlyReg(2);
    rg_man_output[79] = readOnlyReg(3);
    rg_man_output[80] = readOnlyReg(0);
    rg_man_output[81] = readOnlyReg(1);
    rg_man_output[82] = readOnlyReg(2);
    rg_man_output[83] = readOnlyReg(3);
    rg_man_output[84] = readOnlyReg(0);
    rg_man_output[85] = readOnlyReg(1);
    rg_man_output[86] = readOnlyReg(2);
    rg_man_output[87] = readOnlyReg(3);
    rg_man_output[88] = readOnlyReg(0);
    rg_man_output[89] = readOnlyReg(1);
    rg_man_output[90] = readOnlyReg(2);
    rg_man_output[91] = readOnlyReg(3);
    rg_man_output[92] = readOnlyReg(0);
    rg_man_output[93] = readOnlyReg(1);
    rg_man_output[94] = readOnlyReg(2);
    rg_man_output[95] = readOnlyReg(3);
    rg_man_output[96] = readOnlyReg(0);
    rg_man_output[97] = readOnlyReg(1);
    rg_man_output[98] = readOnlyReg(2);
    rg_man_output[99] = readOnlyReg(3);
    rg_man_output[100] = readOnlyReg(0);
    rg_man_output[101] = readOnlyReg(1);
    rg_man_output[102] = readOnlyReg(2);
    rg_man_output[103] = readOnlyReg(3);
    rg_man_output[104] = readOnlyReg(0);
    rg_man_output[105] = readOnlyReg(1);
    rg_man_output[106] = readOnlyReg(2);
    rg_man_output[107] = readOnlyReg(3);
    rg_man_output[108] = readOnlyReg(0);
    rg_man_output[109] = readOnlyReg(1);
    rg_man_output[110] = readOnlyReg(2);
    rg_man_output[111] = readOnlyReg(3);
    rg_man_output[112] = readOnlyReg(0);
    rg_man_output[113] = readOnlyReg(1);
    rg_man_output[114] = readOnlyReg(2);
    rg_man_output[115] = readOnlyReg(3);
    rg_man_output[116] = readOnlyReg(0);
    rg_man_output[117] = readOnlyReg(1);
    rg_man_output[118] = readOnlyReg(2);
    rg_man_output[119] = readOnlyReg(3);
    rg_man_output[120] = readOnlyReg(0);
    rg_man_output[121] = readOnlyReg(1);
    rg_man_output[122] = readOnlyReg(2);
    rg_man_output[123] = readOnlyReg(3);
    rg_man_output[124] = readOnlyReg(0);
    rg_man_output[125] = readOnlyReg(1);
    rg_man_output[126] = readOnlyReg(2);
    rg_man_output[127] = readOnlyReg(3);
    rg_man_output[128] = readOnlyReg(0);
    rg_man_output[129] = readOnlyReg(1);
    rg_man_output[130] = readOnlyReg(2);
    rg_man_output[131] = readOnlyReg(3);
    rg_man_output[132] = readOnlyReg(0);
    rg_man_output[133] = readOnlyReg(1);
    rg_man_output[134] = readOnlyReg(2);
    rg_man_output[135] = readOnlyReg(3);
    rg_man_output[136] = readOnlyReg(0);
    rg_man_output[137] = readOnlyReg(1);
    rg_man_output[138] = readOnlyReg(2);
    rg_man_output[139] = readOnlyReg(3);
    rg_man_output[140] = readOnlyReg(0);
    rg_man_output[141] = readOnlyReg(1);
    rg_man_output[142] = readOnlyReg(2);
    rg_man_output[143] = readOnlyReg(3);
    rg_man_output[144] = readOnlyReg(0);
    rg_man_output[145] = readOnlyReg(1);
    rg_man_output[146] = readOnlyReg(2);
    rg_man_output[147] = readOnlyReg(3);
    rg_man_output[148] = readOnlyReg(0);
    rg_man_output[149] = readOnlyReg(1);
    rg_man_output[150] = readOnlyReg(2);
    rg_man_output[151] = readOnlyReg(3);
    rg_man_output[152] = readOnlyReg(0);
    rg_man_output[153] = readOnlyReg(1);
    rg_man_output[154] = readOnlyReg(2);
    rg_man_output[155] = readOnlyReg(3);
    rg_man_output[156] = readOnlyReg(0);
    rg_man_output[157] = readOnlyReg(1);
    rg_man_output[158] = readOnlyReg(2);
    rg_man_output[159] = readOnlyReg(3);
    rg_man_output[160] = readOnlyReg(0);
    rg_man_output[161] = readOnlyReg(1);
    rg_man_output[162] = readOnlyReg(2);
    rg_man_output[163] = readOnlyReg(3);
    rg_man_output[164] = readOnlyReg(0);
    rg_man_output[165] = readOnlyReg(1);
    rg_man_output[166] = readOnlyReg(2);
    rg_man_output[167] = readOnlyReg(3);
    rg_man_output[168] = readOnlyReg(0);
    rg_man_output[169] = readOnlyReg(1);
    rg_man_output[170] = readOnlyReg(2);
    rg_man_output[171] = readOnlyReg(3);
    rg_man_output[172] = readOnlyReg(0);
    rg_man_output[173] = readOnlyReg(1);
    rg_man_output[174] = readOnlyReg(2);
    rg_man_output[175] = readOnlyReg(3);
    rg_man_output[176] = readOnlyReg(0);
    rg_man_output[177] = readOnlyReg(1);
    rg_man_output[178] = readOnlyReg(2);
    rg_man_output[179] = readOnlyReg(3);
    rg_man_output[180] = readOnlyReg(0);
    rg_man_output[181] = readOnlyReg(1);
    rg_man_output[182] = readOnlyReg(2);
    rg_man_output[183] = readOnlyReg(3);
    rg_man_output[184] = readOnlyReg(0);
    rg_man_output[185] = readOnlyReg(1);
    rg_man_output[186] = readOnlyReg(2);
    rg_man_output[187] = readOnlyReg(3);
    rg_man_output[188] = readOnlyReg(0);
    rg_man_output[189] = readOnlyReg(1);
    rg_man_output[190] = readOnlyReg(2);
    rg_man_output[191] = readOnlyReg(3);
    rg_man_output[192] = readOnlyReg(0);
    rg_man_output[193] = readOnlyReg(1);
    rg_man_output[194] = readOnlyReg(2);
    rg_man_output[195] = readOnlyReg(3);
    rg_man_output[196] = readOnlyReg(0);
    rg_man_output[197] = readOnlyReg(1);
    rg_man_output[198] = readOnlyReg(2);
    rg_man_output[199] = readOnlyReg(3);
    rg_man_output[200] = readOnlyReg(0);
    rg_man_output[201] = readOnlyReg(1);
    rg_man_output[202] = readOnlyReg(2);
    rg_man_output[203] = readOnlyReg(3);
    rg_man_output[204] = readOnlyReg(0);
    rg_man_output[205] = readOnlyReg(1);
    rg_man_output[206] = readOnlyReg(2);
    rg_man_output[207] = readOnlyReg(3);
    rg_man_output[208] = readOnlyReg(0);
    rg_man_output[209] = readOnlyReg(1);
    rg_man_output[210] = readOnlyReg(2);
    rg_man_output[211] = readOnlyReg(3);
    rg_man_output[212] = readOnlyReg(0);
    rg_man_output[213] = readOnlyReg(1);
    rg_man_output[214] = readOnlyReg(2);
    rg_man_output[215] = readOnlyReg(3);
    rg_man_output[216] = readOnlyReg(0);
    rg_man_output[217] = readOnlyReg(1);
    rg_man_output[218] = readOnlyReg(2);
    rg_man_output[219] = readOnlyReg(3);
    rg_man_output[220] = readOnlyReg(0);
    rg_man_output[221] = readOnlyReg(1);
    rg_man_output[222] = readOnlyReg(2);
    rg_man_output[223] = readOnlyReg(3);
    rg_man_output[224] = readOnlyReg(0);
    rg_man_output[225] = readOnlyReg(1);
    rg_man_output[226] = readOnlyReg(2);
    rg_man_output[227] = readOnlyReg(3);
    rg_man_output[228] = readOnlyReg(0);
    rg_man_output[229] = readOnlyReg(1);
    rg_man_output[230] = readOnlyReg(2);
    rg_man_output[231] = readOnlyReg(3);
    rg_man_output[232] = readOnlyReg(0);
    rg_man_output[233] = readOnlyReg(1);
    rg_man_output[234] = readOnlyReg(2);
    rg_man_output[235] = readOnlyReg(3);
    rg_man_output[236] = readOnlyReg(0);
    rg_man_output[237] = readOnlyReg(1);
    rg_man_output[238] = readOnlyReg(2);
    rg_man_output[239] = readOnlyReg(3);
    rg_man_output[240] = readOnlyReg(0);
    rg_man_output[241] = readOnlyReg(1);
    rg_man_output[242] = readOnlyReg(2);
    rg_man_output[243] = readOnlyReg(3);
    rg_man_output[244] = readOnlyReg(0);
    rg_man_output[245] = readOnlyReg(1);
    rg_man_output[246] = readOnlyReg(2);
    rg_man_output[247] = readOnlyReg(3);
    rg_man_output[248] = readOnlyReg(0);
    rg_man_output[249] = readOnlyReg(0);
    rg_man_output[250] = readOnlyReg(0);
    rg_man_output[251] = readOnlyReg(2);
    rg_man_output[252] = readOnlyReg(0);
    rg_man_output[253] = readOnlyReg(1);
    rg_man_output[254] = readOnlyReg(2);
    rg_man_output[255] = readOnlyReg(3);
    rg_man_output[256] = readOnlyReg(0);
    rg_man_output[257] = readOnlyReg(1);
    rg_man_output[258] = readOnlyReg(2);
    rg_man_output[259] = readOnlyReg(3);
    rg_man_output[260] = readOnlyReg(0);
    rg_man_output[261] = readOnlyReg(1);
    rg_man_output[262] = readOnlyReg(2);
    rg_man_output[263] = readOnlyReg(3);
    rg_man_output[264] = readOnlyReg(0);
    rg_man_output[265] = readOnlyReg(1);
    rg_man_output[266] = readOnlyReg(2);
    rg_man_output[267] = readOnlyReg(3);
    rg_man_output[268] = readOnlyReg(0);
    rg_man_output[269] = readOnlyReg(1);
    rg_man_output[270] = readOnlyReg(2);
    rg_man_output[271] = readOnlyReg(3);
    rg_man_output[272] = readOnlyReg(0);
    rg_man_output[273] = readOnlyReg(1);
    rg_man_output[274] = readOnlyReg(2);
    rg_man_output[275] = readOnlyReg(3);
    rg_man_output[276] = readOnlyReg(0);
    rg_man_output[277] = readOnlyReg(1);
    rg_man_output[278] = readOnlyReg(2);
    rg_man_output[279] = readOnlyReg(3);
    rg_man_output[280] = readOnlyReg(0);
    rg_man_output[281] = readOnlyReg(1);
    rg_man_output[282] = readOnlyReg(2);
    rg_man_output[283] = readOnlyReg(3);
    rg_man_output[284] = readOnlyReg(0);
    rg_man_output[285] = readOnlyReg(1);
    rg_man_output[286] = readOnlyReg(2);
    rg_man_output[287] = readOnlyReg(3);
    rg_man_output[288] = readOnlyReg(0);
    rg_man_output[289] = readOnlyReg(1);
    rg_man_output[290] = readOnlyReg(2);
    rg_man_output[291] = readOnlyReg(3);
    rg_man_output[292] = readOnlyReg(0);
    rg_man_output[293] = readOnlyReg(1);
    rg_man_output[294] = readOnlyReg(2);
    rg_man_output[295] = readOnlyReg(3);
    rg_man_output[296] = readOnlyReg(0);
    rg_man_output[297] = readOnlyReg(1);
    rg_man_output[298] = readOnlyReg(2);
    rg_man_output[299] = readOnlyReg(3);
    rg_man_output[300] = readOnlyReg(0);
    rg_man_output[301] = readOnlyReg(1);
    rg_man_output[302] = readOnlyReg(2);
    rg_man_output[303] = readOnlyReg(3);
    rg_man_output[304] = readOnlyReg(0);
    rg_man_output[305] = readOnlyReg(1);
    rg_man_output[306] = readOnlyReg(2);
    rg_man_output[307] = readOnlyReg(3);
    rg_man_output[308] = readOnlyReg(0);
    rg_man_output[309] = readOnlyReg(1);
    rg_man_output[310] = readOnlyReg(2);
    rg_man_output[311] = readOnlyReg(3);
    rg_man_output[312] = readOnlyReg(0);
    rg_man_output[313] = readOnlyReg(1);
    rg_man_output[314] = readOnlyReg(2);
    rg_man_output[315] = readOnlyReg(3);
    rg_man_output[316] = readOnlyReg(0);
    rg_man_output[317] = readOnlyReg(1);
    rg_man_output[318] = readOnlyReg(2);
    rg_man_output[319] = readOnlyReg(3);
    rg_man_output[320] = readOnlyReg(0);
    rg_man_output[321] = readOnlyReg(1);
    rg_man_output[322] = readOnlyReg(2);
    rg_man_output[323] = readOnlyReg(3);
    rg_man_output[324] = readOnlyReg(0);
    rg_man_output[325] = readOnlyReg(1);
    rg_man_output[326] = readOnlyReg(2);
    rg_man_output[327] = readOnlyReg(3);
    rg_man_output[328] = readOnlyReg(0);
    rg_man_output[329] = readOnlyReg(1);
    rg_man_output[330] = readOnlyReg(2);
    rg_man_output[331] = readOnlyReg(3);
    rg_man_output[332] = readOnlyReg(0);
    rg_man_output[333] = readOnlyReg(1);
    rg_man_output[334] = readOnlyReg(2);
    rg_man_output[335] = readOnlyReg(3);
    rg_man_output[336] = readOnlyReg(0);
    rg_man_output[337] = readOnlyReg(1);
    rg_man_output[338] = readOnlyReg(2);
    rg_man_output[339] = readOnlyReg(3);
    rg_man_output[340] = readOnlyReg(0);
    rg_man_output[341] = readOnlyReg(1);
    rg_man_output[342] = readOnlyReg(2);
    rg_man_output[343] = readOnlyReg(3);
    rg_man_output[344] = readOnlyReg(0);
    rg_man_output[345] = readOnlyReg(1);
    rg_man_output[346] = readOnlyReg(2);
    rg_man_output[347] = readOnlyReg(3);
    rg_man_output[348] = readOnlyReg(0);
    rg_man_output[349] = readOnlyReg(1);
    rg_man_output[350] = readOnlyReg(2);
    rg_man_output[351] = readOnlyReg(3);
    rg_man_output[352] = readOnlyReg(0);
    rg_man_output[353] = readOnlyReg(1);
    rg_man_output[354] = readOnlyReg(2);
    rg_man_output[355] = readOnlyReg(3);
    rg_man_output[356] = readOnlyReg(0);
    rg_man_output[357] = readOnlyReg(1);
    rg_man_output[358] = readOnlyReg(2);
    rg_man_output[359] = readOnlyReg(3);
    rg_man_output[360] = readOnlyReg(0);
    rg_man_output[361] = readOnlyReg(1);
    rg_man_output[362] = readOnlyReg(2);
    rg_man_output[363] = readOnlyReg(3);
    rg_man_output[364] = readOnlyReg(0);
    rg_man_output[365] = readOnlyReg(1);
    rg_man_output[366] = readOnlyReg(2);
    rg_man_output[367] = readOnlyReg(3);
    rg_man_output[368] = readOnlyReg(0);
    rg_man_output[369] = readOnlyReg(1);
    rg_man_output[370] = readOnlyReg(2);
    rg_man_output[371] = readOnlyReg(3);
    rg_man_output[372] = readOnlyReg(0);
    rg_man_output[373] = readOnlyReg(1);
    rg_man_output[374] = readOnlyReg(2);
    rg_man_output[375] = readOnlyReg(3);

    Reg#(Int#(5)) rg_exp_output[376];
    rg_exp_output[0] = readOnlyReg(-62);
    rg_exp_output[1] = readOnlyReg(-62);
    rg_exp_output[2] = readOnlyReg(-62);
    rg_exp_output[3] = readOnlyReg(-62);
    rg_exp_output[4] = readOnlyReg(-61);
    rg_exp_output[5] = readOnlyReg(-61);
    rg_exp_output[6] = readOnlyReg(-61);
    rg_exp_output[7] = readOnlyReg(-61);
    rg_exp_output[8] = readOnlyReg(-60);
    rg_exp_output[9] = readOnlyReg(-60);
    rg_exp_output[10] = readOnlyReg(-60);
    rg_exp_output[11] = readOnlyReg(-60);
    rg_exp_output[12] = readOnlyReg(-59);
    rg_exp_output[13] = readOnlyReg(-59);
    rg_exp_output[14] = readOnlyReg(-59);
    rg_exp_output[15] = readOnlyReg(-59);
    rg_exp_output[16] = readOnlyReg(-58);
    rg_exp_output[17] = readOnlyReg(-58);
    rg_exp_output[18] = readOnlyReg(-58);
    rg_exp_output[19] = readOnlyReg(-58);
    rg_exp_output[20] = readOnlyReg(-57);
    rg_exp_output[21] = readOnlyReg(-57);
    rg_exp_output[22] = readOnlyReg(-57);
    rg_exp_output[23] = readOnlyReg(-57);
    rg_exp_output[24] = readOnlyReg(-56);
    rg_exp_output[25] = readOnlyReg(-56);
    rg_exp_output[26] = readOnlyReg(-56);
    rg_exp_output[27] = readOnlyReg(-56);
    rg_exp_output[28] = readOnlyReg(-55);
    rg_exp_output[29] = readOnlyReg(-55);
    rg_exp_output[30] = readOnlyReg(-55);
    rg_exp_output[31] = readOnlyReg(-55);
    rg_exp_output[32] = readOnlyReg(-54);
    rg_exp_output[33] = readOnlyReg(-54);
    rg_exp_output[34] = readOnlyReg(-54);
    rg_exp_output[35] = readOnlyReg(-54);
    rg_exp_output[36] = readOnlyReg(-53);
    rg_exp_output[37] = readOnlyReg(-53);
    rg_exp_output[38] = readOnlyReg(-53);
    rg_exp_output[39] = readOnlyReg(-53);
    rg_exp_output[40] = readOnlyReg(-52);
    rg_exp_output[41] = readOnlyReg(-52);
    rg_exp_output[42] = readOnlyReg(-52);
    rg_exp_output[43] = readOnlyReg(-52);
    rg_exp_output[44] = readOnlyReg(-51);
    rg_exp_output[45] = readOnlyReg(-51);
    rg_exp_output[46] = readOnlyReg(-51);
    rg_exp_output[47] = readOnlyReg(-51);
    rg_exp_output[48] = readOnlyReg(-50);
    rg_exp_output[49] = readOnlyReg(-50);
    rg_exp_output[50] = readOnlyReg(-50);
    rg_exp_output[51] = readOnlyReg(-50);
    rg_exp_output[52] = readOnlyReg(-49);
    rg_exp_output[53] = readOnlyReg(-49);
    rg_exp_output[54] = readOnlyReg(-49);
    rg_exp_output[55] = readOnlyReg(-49);
    rg_exp_output[56] = readOnlyReg(-48);
    rg_exp_output[57] = readOnlyReg(-48);
    rg_exp_output[58] = readOnlyReg(-48);
    rg_exp_output[59] = readOnlyReg(-48);
    rg_exp_output[60] = readOnlyReg(-47);
    rg_exp_output[61] = readOnlyReg(-47);
    rg_exp_output[62] = readOnlyReg(-47);
    rg_exp_output[63] = readOnlyReg(-47);
    rg_exp_output[64] = readOnlyReg(-46);
    rg_exp_output[65] = readOnlyReg(-46);
    rg_exp_output[66] = readOnlyReg(-46);
    rg_exp_output[67] = readOnlyReg(-46);
    rg_exp_output[68] = readOnlyReg(-45);
    rg_exp_output[69] = readOnlyReg(-45);
    rg_exp_output[70] = readOnlyReg(-45);
    rg_exp_output[71] = readOnlyReg(-45);
    rg_exp_output[72] = readOnlyReg(-44);
    rg_exp_output[73] = readOnlyReg(-44);
    rg_exp_output[74] = readOnlyReg(-44);
    rg_exp_output[75] = readOnlyReg(-44);
    rg_exp_output[76] = readOnlyReg(-43);
    rg_exp_output[77] = readOnlyReg(-43);
    rg_exp_output[78] = readOnlyReg(-43);
    rg_exp_output[79] = readOnlyReg(-43);
    rg_exp_output[80] = readOnlyReg(-42);
    rg_exp_output[81] = readOnlyReg(-42);
    rg_exp_output[82] = readOnlyReg(-42);
    rg_exp_output[83] = readOnlyReg(-42);
    rg_exp_output[84] = readOnlyReg(-41);
    rg_exp_output[85] = readOnlyReg(-41);
    rg_exp_output[86] = readOnlyReg(-41);
    rg_exp_output[87] = readOnlyReg(-41);
    rg_exp_output[88] = readOnlyReg(-40);
    rg_exp_output[89] = readOnlyReg(-40);
    rg_exp_output[90] = readOnlyReg(-40);
    rg_exp_output[91] = readOnlyReg(-40);
    rg_exp_output[92] = readOnlyReg(-39);
    rg_exp_output[93] = readOnlyReg(-39);
    rg_exp_output[94] = readOnlyReg(-39);
    rg_exp_output[95] = readOnlyReg(-39);
    rg_exp_output[96] = readOnlyReg(-38);
    rg_exp_output[97] = readOnlyReg(-38);
    rg_exp_output[98] = readOnlyReg(-38);
    rg_exp_output[99] = readOnlyReg(-38);
    rg_exp_output[100] = readOnlyReg(-37);
    rg_exp_output[101] = readOnlyReg(-37);
    rg_exp_output[102] = readOnlyReg(-37);
    rg_exp_output[103] = readOnlyReg(-37);
    rg_exp_output[104] = readOnlyReg(-36);
    rg_exp_output[105] = readOnlyReg(-36);
    rg_exp_output[106] = readOnlyReg(-36);
    rg_exp_output[107] = readOnlyReg(-36);
    rg_exp_output[108] = readOnlyReg(-35);
    rg_exp_output[109] = readOnlyReg(-35);
    rg_exp_output[110] = readOnlyReg(-35);
    rg_exp_output[111] = readOnlyReg(-35);
    rg_exp_output[112] = readOnlyReg(-34);
    rg_exp_output[113] = readOnlyReg(-34);
    rg_exp_output[114] = readOnlyReg(-34);
    rg_exp_output[115] = readOnlyReg(-34);
    rg_exp_output[116] = readOnlyReg(-33);
    rg_exp_output[117] = readOnlyReg(-33);
    rg_exp_output[118] = readOnlyReg(-33);
    rg_exp_output[119] = readOnlyReg(-33);
    rg_exp_output[120] = readOnlyReg(-32);
    rg_exp_output[121] = readOnlyReg(-32);
    rg_exp_output[122] = readOnlyReg(-32);
    rg_exp_output[123] = readOnlyReg(-32);
    rg_exp_output[124] = readOnlyReg(-31);
    rg_exp_output[125] = readOnlyReg(-31);
    rg_exp_output[126] = readOnlyReg(-31);
    rg_exp_output[127] = readOnlyReg(-31);
    rg_exp_output[128] = readOnlyReg(-30);
    rg_exp_output[129] = readOnlyReg(-30);
    rg_exp_output[130] = readOnlyReg(-30);
    rg_exp_output[131] = readOnlyReg(-30);
    rg_exp_output[132] = readOnlyReg(-29);
    rg_exp_output[133] = readOnlyReg(-29);
    rg_exp_output[134] = readOnlyReg(-29);
    rg_exp_output[135] = readOnlyReg(-29);
    rg_exp_output[136] = readOnlyReg(-28);
    rg_exp_output[137] = readOnlyReg(-28);
    rg_exp_output[138] = readOnlyReg(-28);
    rg_exp_output[139] = readOnlyReg(-28);
    rg_exp_output[140] = readOnlyReg(-27);
    rg_exp_output[141] = readOnlyReg(-27);
    rg_exp_output[142] = readOnlyReg(-27);
    rg_exp_output[143] = readOnlyReg(-27);
    rg_exp_output[144] = readOnlyReg(-26);
    rg_exp_output[145] = readOnlyReg(-26);
    rg_exp_output[146] = readOnlyReg(-26);
    rg_exp_output[147] = readOnlyReg(-26);
    rg_exp_output[148] = readOnlyReg(-25);
    rg_exp_output[149] = readOnlyReg(-25);
    rg_exp_output[150] = readOnlyReg(-25);
    rg_exp_output[151] = readOnlyReg(-25);
    rg_exp_output[152] = readOnlyReg(-24);
    rg_exp_output[153] = readOnlyReg(-24);
    rg_exp_output[154] = readOnlyReg(-24);
    rg_exp_output[155] = readOnlyReg(-24);
    rg_exp_output[156] = readOnlyReg(-23);
    rg_exp_output[157] = readOnlyReg(-23);
    rg_exp_output[158] = readOnlyReg(-23);
    rg_exp_output[159] = readOnlyReg(-23);
    rg_exp_output[160] = readOnlyReg(-22);
    rg_exp_output[161] = readOnlyReg(-22);
    rg_exp_output[162] = readOnlyReg(-22);
    rg_exp_output[163] = readOnlyReg(-22);
    rg_exp_output[164] = readOnlyReg(-21);
    rg_exp_output[165] = readOnlyReg(-21);
    rg_exp_output[166] = readOnlyReg(-21);
    rg_exp_output[167] = readOnlyReg(-21);
    rg_exp_output[168] = readOnlyReg(-20);
    rg_exp_output[169] = readOnlyReg(-20);
    rg_exp_output[170] = readOnlyReg(-20);
    rg_exp_output[171] = readOnlyReg(-20);
    rg_exp_output[172] = readOnlyReg(-19);
    rg_exp_output[173] = readOnlyReg(-19);
    rg_exp_output[174] = readOnlyReg(-19);
    rg_exp_output[175] = readOnlyReg(-19);
    rg_exp_output[176] = readOnlyReg(-18);
    rg_exp_output[177] = readOnlyReg(-18);
    rg_exp_output[178] = readOnlyReg(-18);
    rg_exp_output[179] = readOnlyReg(-18);
    rg_exp_output[180] = readOnlyReg(-17);
    rg_exp_output[181] = readOnlyReg(-17);
    rg_exp_output[182] = readOnlyReg(-17);
    rg_exp_output[183] = readOnlyReg(-17);
    rg_exp_output[184] = readOnlyReg(-16);
    rg_exp_output[185] = readOnlyReg(-16);
    rg_exp_output[186] = readOnlyReg(-16);
    rg_exp_output[187] = readOnlyReg(-16);
    rg_exp_output[188] = readOnlyReg(-15);
    rg_exp_output[189] = readOnlyReg(-15);
    rg_exp_output[190] = readOnlyReg(-15);
    rg_exp_output[191] = readOnlyReg(-15);
    rg_exp_output[192] = readOnlyReg(-14);
    rg_exp_output[193] = readOnlyReg(-14);
    rg_exp_output[194] = readOnlyReg(-14);
    rg_exp_output[195] = readOnlyReg(-14);
    rg_exp_output[196] = readOnlyReg(-13);
    rg_exp_output[197] = readOnlyReg(-13);
    rg_exp_output[198] = readOnlyReg(-13);
    rg_exp_output[199] = readOnlyReg(-13);
    rg_exp_output[200] = readOnlyReg(-12);
    rg_exp_output[201] = readOnlyReg(-12);
    rg_exp_output[202] = readOnlyReg(-12);
    rg_exp_output[203] = readOnlyReg(-12);
    rg_exp_output[204] = readOnlyReg(-11);
    rg_exp_output[205] = readOnlyReg(-11);
    rg_exp_output[206] = readOnlyReg(-11);
    rg_exp_output[207] = readOnlyReg(-11);
    rg_exp_output[208] = readOnlyReg(-10);
    rg_exp_output[209] = readOnlyReg(-10);
    rg_exp_output[210] = readOnlyReg(-10);
    rg_exp_output[211] = readOnlyReg(-10);
    rg_exp_output[212] = readOnlyReg(-9);
    rg_exp_output[213] = readOnlyReg(-9);
    rg_exp_output[214] = readOnlyReg(-9);
    rg_exp_output[215] = readOnlyReg(-9);
    rg_exp_output[216] = readOnlyReg(-8);
    rg_exp_output[217] = readOnlyReg(-8);
    rg_exp_output[218] = readOnlyReg(-8);
    rg_exp_output[219] = readOnlyReg(-8);
    rg_exp_output[220] = readOnlyReg(-7);
    rg_exp_output[221] = readOnlyReg(-7);
    rg_exp_output[222] = readOnlyReg(-7);
    rg_exp_output[223] = readOnlyReg(-7);
    rg_exp_output[224] = readOnlyReg(-6);
    rg_exp_output[225] = readOnlyReg(-6);
    rg_exp_output[226] = readOnlyReg(-6);
    rg_exp_output[227] = readOnlyReg(-6);
    rg_exp_output[228] = readOnlyReg(-5);
    rg_exp_output[229] = readOnlyReg(-5);
    rg_exp_output[230] = readOnlyReg(-5);
    rg_exp_output[231] = readOnlyReg(-5);
    rg_exp_output[232] = readOnlyReg(-4);
    rg_exp_output[233] = readOnlyReg(-4);
    rg_exp_output[234] = readOnlyReg(-4);
    rg_exp_output[235] = readOnlyReg(-4);
    rg_exp_output[236] = readOnlyReg(-3);
    rg_exp_output[237] = readOnlyReg(-3);
    rg_exp_output[238] = readOnlyReg(-3);
    rg_exp_output[239] = readOnlyReg(-3);
    rg_exp_output[240] = readOnlyReg(-2);
    rg_exp_output[241] = readOnlyReg(-2);
    rg_exp_output[242] = readOnlyReg(-2);
    rg_exp_output[243] = readOnlyReg(-2);
    rg_exp_output[244] = readOnlyReg(-1);
    rg_exp_output[245] = readOnlyReg(-1);
    rg_exp_output[246] = readOnlyReg(-1);
    rg_exp_output[247] = readOnlyReg(-1);
    rg_exp_output[248] = readOnlyReg(0);
    rg_exp_output[249] = readOnlyReg(-2);
    rg_exp_output[250] = readOnlyReg(-1);
    rg_exp_output[251] = readOnlyReg(-1);
    rg_exp_output[252] = readOnlyReg(1);
    rg_exp_output[253] = readOnlyReg(1);
    rg_exp_output[254] = readOnlyReg(1);
    rg_exp_output[255] = readOnlyReg(1);
    rg_exp_output[256] = readOnlyReg(2);
    rg_exp_output[257] = readOnlyReg(2);
    rg_exp_output[258] = readOnlyReg(2);
    rg_exp_output[259] = readOnlyReg(2);
    rg_exp_output[260] = readOnlyReg(3);
    rg_exp_output[261] = readOnlyReg(3);
    rg_exp_output[262] = readOnlyReg(3);
    rg_exp_output[263] = readOnlyReg(3);
    rg_exp_output[264] = readOnlyReg(4);
    rg_exp_output[265] = readOnlyReg(4);
    rg_exp_output[266] = readOnlyReg(4);
    rg_exp_output[267] = readOnlyReg(4);
    rg_exp_output[268] = readOnlyReg(5);
    rg_exp_output[269] = readOnlyReg(5);
    rg_exp_output[270] = readOnlyReg(5);
    rg_exp_output[271] = readOnlyReg(5);
    rg_exp_output[272] = readOnlyReg(6);
    rg_exp_output[273] = readOnlyReg(6);
    rg_exp_output[274] = readOnlyReg(6);
    rg_exp_output[275] = readOnlyReg(6);
    rg_exp_output[276] = readOnlyReg(7);
    rg_exp_output[277] = readOnlyReg(7);
    rg_exp_output[278] = readOnlyReg(7);
    rg_exp_output[279] = readOnlyReg(7);
    rg_exp_output[280] = readOnlyReg(8);
    rg_exp_output[281] = readOnlyReg(8);
    rg_exp_output[282] = readOnlyReg(8);
    rg_exp_output[283] = readOnlyReg(8);
    rg_exp_output[284] = readOnlyReg(9);
    rg_exp_output[285] = readOnlyReg(9);
    rg_exp_output[286] = readOnlyReg(9);
    rg_exp_output[287] = readOnlyReg(9);
    rg_exp_output[288] = readOnlyReg(10);
    rg_exp_output[289] = readOnlyReg(10);
    rg_exp_output[290] = readOnlyReg(10);
    rg_exp_output[291] = readOnlyReg(10);
    rg_exp_output[292] = readOnlyReg(11);
    rg_exp_output[293] = readOnlyReg(11);
    rg_exp_output[294] = readOnlyReg(11);
    rg_exp_output[295] = readOnlyReg(11);
    rg_exp_output[296] = readOnlyReg(12);
    rg_exp_output[297] = readOnlyReg(12);
    rg_exp_output[298] = readOnlyReg(12);
    rg_exp_output[299] = readOnlyReg(12);
    rg_exp_output[300] = readOnlyReg(13);
    rg_exp_output[301] = readOnlyReg(13);
    rg_exp_output[302] = readOnlyReg(13);
    rg_exp_output[303] = readOnlyReg(13);
    rg_exp_output[304] = readOnlyReg(14);
    rg_exp_output[305] = readOnlyReg(14);
    rg_exp_output[306] = readOnlyReg(14);
    rg_exp_output[307] = readOnlyReg(14);
    rg_exp_output[308] = readOnlyReg(15);
    rg_exp_output[309] = readOnlyReg(15);
    rg_exp_output[310] = readOnlyReg(15);
    rg_exp_output[311] = readOnlyReg(15);
    rg_exp_output[312] = readOnlyReg(16);
    rg_exp_output[313] = readOnlyReg(16);
    rg_exp_output[314] = readOnlyReg(16);
    rg_exp_output[315] = readOnlyReg(16);
    rg_exp_output[316] = readOnlyReg(17);
    rg_exp_output[317] = readOnlyReg(17);
    rg_exp_output[318] = readOnlyReg(17);
    rg_exp_output[319] = readOnlyReg(17);
    rg_exp_output[320] = readOnlyReg(18);
    rg_exp_output[321] = readOnlyReg(18);
    rg_exp_output[322] = readOnlyReg(18);
    rg_exp_output[323] = readOnlyReg(18);
    rg_exp_output[324] = readOnlyReg(19);
    rg_exp_output[325] = readOnlyReg(19);
    rg_exp_output[326] = readOnlyReg(19);
    rg_exp_output[327] = readOnlyReg(19);
    rg_exp_output[328] = readOnlyReg(20);
    rg_exp_output[329] = readOnlyReg(20);
    rg_exp_output[330] = readOnlyReg(20);
    rg_exp_output[331] = readOnlyReg(20);
    rg_exp_output[332] = readOnlyReg(21);
    rg_exp_output[333] = readOnlyReg(21);
    rg_exp_output[334] = readOnlyReg(21);
    rg_exp_output[335] = readOnlyReg(21);
    rg_exp_output[336] = readOnlyReg(22);
    rg_exp_output[337] = readOnlyReg(22);
    rg_exp_output[338] = readOnlyReg(22);
    rg_exp_output[339] = readOnlyReg(22);
    rg_exp_output[340] = readOnlyReg(23);
    rg_exp_output[341] = readOnlyReg(23);
    rg_exp_output[342] = readOnlyReg(23);
    rg_exp_output[343] = readOnlyReg(23);
    rg_exp_output[344] = readOnlyReg(24);
    rg_exp_output[345] = readOnlyReg(24);
    rg_exp_output[346] = readOnlyReg(24);
    rg_exp_output[347] = readOnlyReg(24);
    rg_exp_output[348] = readOnlyReg(25);
    rg_exp_output[349] = readOnlyReg(25);
    rg_exp_output[350] = readOnlyReg(25);
    rg_exp_output[351] = readOnlyReg(25);
    rg_exp_output[352] = readOnlyReg(26);
    rg_exp_output[353] = readOnlyReg(26);
    rg_exp_output[354] = readOnlyReg(26);
    rg_exp_output[355] = readOnlyReg(26);
    rg_exp_output[356] = readOnlyReg(27);
    rg_exp_output[357] = readOnlyReg(27);
    rg_exp_output[358] = readOnlyReg(27);
    rg_exp_output[359] = readOnlyReg(27);
    rg_exp_output[360] = readOnlyReg(28);
    rg_exp_output[361] = readOnlyReg(28);
    rg_exp_output[362] = readOnlyReg(28);
    rg_exp_output[363] = readOnlyReg(28);
    rg_exp_output[364] = readOnlyReg(29);
    rg_exp_output[365] = readOnlyReg(29);
    rg_exp_output[366] = readOnlyReg(29);
    rg_exp_output[367] = readOnlyReg(29);
    rg_exp_output[368] = readOnlyReg(30);
    rg_exp_output[369] = readOnlyReg(30);
    rg_exp_output[370] = readOnlyReg(30);
    rg_exp_output[371] = readOnlyReg(30);
    rg_exp_output[372] = readOnlyReg(31);
    rg_exp_output[373] = readOnlyReg(31);
    rg_exp_output[374] = readOnlyReg(31);
    rg_exp_output[375] = readOnlyReg(31);

    method Tuple2#(Bit#(5), Bit#(2)) mv_sig_output(Bit#(4) exp, Bit#(2) man);
      Bit#(6) index = {man, exp};
      return tuple2(rg_man_output[index], rg_exp_output[index]);
    endmethod
  endmodule

  interface Ifc_sigmoid_lut_region_3;
    method Tuple2#(Int#(7), Bit#(2)) mv_sig_output(Bit#(2) exp, Bit#(2) man);
  endinterface

  module mksigmoid_lut_region_3(Ifc_sigmoid_lut_region_3);
    Reg#(Bit#(2)) rg_man_output[350];
    rg_man_output[0] = readOnlyReg(3);
    rg_man_output[1] = readOnlyReg(3);
    rg_man_output[2] = readOnlyReg(3);
    rg_man_output[3] = readOnlyReg(3);
    rg_man_output[4] = readOnlyReg(1);
    rg_man_output[5] = readOnlyReg(3);
    rg_man_output[6] = readOnlyReg(3);
    rg_man_output[7] = readOnlyReg(1);
    rg_man_output[8] = readOnlyReg(3);
    rg_man_output[9] = readOnlyReg(3);
    rg_man_output[10] = readOnlyReg(1);
    rg_man_output[11] = readOnlyReg(3);
    rg_man_output[12] = readOnlyReg(3);
    rg_man_output[13] = readOnlyReg(1);
    rg_man_output[14] = readOnlyReg(3);
    rg_man_output[15] = readOnlyReg(3);
    rg_man_output[16] = readOnlyReg(1);
    rg_man_output[17] = readOnlyReg(3);
    rg_man_output[18] = readOnlyReg(3);
    rg_man_output[19] = readOnlyReg(1);
    rg_man_output[20] = readOnlyReg(3);
    rg_man_output[21] = readOnlyReg(3);
    rg_man_output[22] = readOnlyReg(1);
    rg_man_output[23] = readOnlyReg(3);
    rg_man_output[24] = readOnlyReg(3);
    rg_man_output[25] = readOnlyReg(1);
    rg_man_output[26] = readOnlyReg(3);
    rg_man_output[27] = readOnlyReg(3);
    rg_man_output[28] = readOnlyReg(1);
    rg_man_output[29] = readOnlyReg(3);
    rg_man_output[30] = readOnlyReg(3);
    rg_man_output[31] = readOnlyReg(1);
    rg_man_output[32] = readOnlyReg(3);
    rg_man_output[33] = readOnlyReg(3);
    rg_man_output[34] = readOnlyReg(1);
    rg_man_output[35] = readOnlyReg(3);
    rg_man_output[36] = readOnlyReg(3);
    rg_man_output[37] = readOnlyReg(1);
    rg_man_output[38] = readOnlyReg(3);
    rg_man_output[39] = readOnlyReg(3);
    rg_man_output[40] = readOnlyReg(1);
    rg_man_output[41] = readOnlyReg(3);
    rg_man_output[42] = readOnlyReg(3);
    rg_man_output[43] = readOnlyReg(1);
    rg_man_output[44] = readOnlyReg(3);
    rg_man_output[45] = readOnlyReg(3);
    rg_man_output[46] = readOnlyReg(1);
    rg_man_output[47] = readOnlyReg(3);
    rg_man_output[48] = readOnlyReg(3);
    rg_man_output[49] = readOnlyReg(1);
    rg_man_output[50] = readOnlyReg(3);
    rg_man_output[51] = readOnlyReg(3);
    rg_man_output[52] = readOnlyReg(1);
    rg_man_output[53] = readOnlyReg(3);
    rg_man_output[54] = readOnlyReg(3);
    rg_man_output[55] = readOnlyReg(1);
    rg_man_output[56] = readOnlyReg(3);
    rg_man_output[57] = readOnlyReg(3);
    rg_man_output[58] = readOnlyReg(1);
    rg_man_output[59] = readOnlyReg(3);
    rg_man_output[60] = readOnlyReg(3);
    rg_man_output[61] = readOnlyReg(1);
    rg_man_output[62] = readOnlyReg(3);
    rg_man_output[63] = readOnlyReg(3);
    rg_man_output[64] = readOnlyReg(1);
    rg_man_output[65] = readOnlyReg(3);
    rg_man_output[66] = readOnlyReg(3);
    rg_man_output[67] = readOnlyReg(1);
    rg_man_output[68] = readOnlyReg(3);
    rg_man_output[69] = readOnlyReg(3);
    rg_man_output[70] = readOnlyReg(1);
    rg_man_output[71] = readOnlyReg(3);
    rg_man_output[72] = readOnlyReg(3);
    rg_man_output[73] = readOnlyReg(1);
    rg_man_output[74] = readOnlyReg(3);
    rg_man_output[75] = readOnlyReg(3);
    rg_man_output[76] = readOnlyReg(1);
    rg_man_output[77] = readOnlyReg(3);
    rg_man_output[78] = readOnlyReg(3);
    rg_man_output[79] = readOnlyReg(1);
    rg_man_output[80] = readOnlyReg(3);
    rg_man_output[81] = readOnlyReg(3);
    rg_man_output[82] = readOnlyReg(1);
    rg_man_output[83] = readOnlyReg(3);
    rg_man_output[84] = readOnlyReg(3);
    rg_man_output[85] = readOnlyReg(1);
    rg_man_output[86] = readOnlyReg(3);
    rg_man_output[87] = readOnlyReg(3);
    rg_man_output[88] = readOnlyReg(1);
    rg_man_output[89] = readOnlyReg(3);
    rg_man_output[90] = readOnlyReg(3);
    rg_man_output[91] = readOnlyReg(1);
    rg_man_output[92] = readOnlyReg(3);
    rg_man_output[93] = readOnlyReg(3);
    rg_man_output[94] = readOnlyReg(1);
    rg_man_output[95] = readOnlyReg(3);
    rg_man_output[96] = readOnlyReg(3);
    rg_man_output[97] = readOnlyReg(1);
    rg_man_output[98] = readOnlyReg(3);
    rg_man_output[99] = readOnlyReg(3);
    rg_man_output[100] = readOnlyReg(1);
    rg_man_output[101] = readOnlyReg(3);
    rg_man_output[102] = readOnlyReg(3);
    rg_man_output[103] = readOnlyReg(1);
    rg_man_output[104] = readOnlyReg(3);
    rg_man_output[105] = readOnlyReg(3);
    rg_man_output[106] = readOnlyReg(1);
    rg_man_output[107] = readOnlyReg(3);
    rg_man_output[108] = readOnlyReg(3);
    rg_man_output[109] = readOnlyReg(1);
    rg_man_output[110] = readOnlyReg(3);
    rg_man_output[111] = readOnlyReg(3);
    rg_man_output[112] = readOnlyReg(1);
    rg_man_output[113] = readOnlyReg(3);
    rg_man_output[114] = readOnlyReg(3);
    rg_man_output[115] = readOnlyReg(1);
    rg_man_output[116] = readOnlyReg(3);
    rg_man_output[117] = readOnlyReg(3);
    rg_man_output[118] = readOnlyReg(1);
    rg_man_output[119] = readOnlyReg(3);
    rg_man_output[120] = readOnlyReg(3);
    rg_man_output[121] = readOnlyReg(1);
    rg_man_output[122] = readOnlyReg(3);
    rg_man_output[123] = readOnlyReg(3);
    rg_man_output[124] = readOnlyReg(1);
    rg_man_output[125] = readOnlyReg(3);
    rg_man_output[126] = readOnlyReg(3);
    rg_man_output[127] = readOnlyReg(1);
    rg_man_output[128] = readOnlyReg(3);
    rg_man_output[129] = readOnlyReg(3);
    rg_man_output[130] = readOnlyReg(1);
    rg_man_output[131] = readOnlyReg(3);
    rg_man_output[132] = readOnlyReg(3);
    rg_man_output[133] = readOnlyReg(1);
    rg_man_output[134] = readOnlyReg(3);
    rg_man_output[135] = readOnlyReg(3);
    rg_man_output[136] = readOnlyReg(1);
    rg_man_output[137] = readOnlyReg(3);
    rg_man_output[138] = readOnlyReg(3);
    rg_man_output[139] = readOnlyReg(1);
    rg_man_output[140] = readOnlyReg(3);
    rg_man_output[141] = readOnlyReg(3);
    rg_man_output[142] = readOnlyReg(1);
    rg_man_output[143] = readOnlyReg(3);
    rg_man_output[144] = readOnlyReg(3);
    rg_man_output[145] = readOnlyReg(1);
    rg_man_output[146] = readOnlyReg(3);
    rg_man_output[147] = readOnlyReg(3);
    rg_man_output[148] = readOnlyReg(1);
    rg_man_output[149] = readOnlyReg(3);
    rg_man_output[150] = readOnlyReg(3);
    rg_man_output[151] = readOnlyReg(1);
    rg_man_output[152] = readOnlyReg(3);
    rg_man_output[153] = readOnlyReg(2);
    rg_man_output[154] = readOnlyReg(0);
    rg_man_output[155] = readOnlyReg(2);
    rg_man_output[156] = readOnlyReg(2);
    rg_man_output[157] = readOnlyReg(3);
    rg_man_output[158] = readOnlyReg(0);
    rg_man_output[159] = readOnlyReg(0);
    rg_man_output[160] = readOnlyReg(0);
    rg_man_output[161] = readOnlyReg(0);
    rg_man_output[162] = readOnlyReg(0);
    rg_man_output[163] = readOnlyReg(0);
    rg_man_output[164] = readOnlyReg(0);
    rg_man_output[165] = readOnlyReg(0);
    rg_man_output[166] = readOnlyReg(2);
    rg_man_output[167] = readOnlyReg(0);
    rg_man_output[168] = readOnlyReg(0);
    rg_man_output[169] = readOnlyReg(2);
    rg_man_output[170] = readOnlyReg(0);
    rg_man_output[171] = readOnlyReg(0);
    rg_man_output[172] = readOnlyReg(2);
    rg_man_output[173] = readOnlyReg(0);
    rg_man_output[174] = readOnlyReg(0);
    rg_man_output[175] = readOnlyReg(2);
    rg_man_output[176] = readOnlyReg(0);
    rg_man_output[177] = readOnlyReg(0);
    rg_man_output[178] = readOnlyReg(2);
    rg_man_output[179] = readOnlyReg(0);
    rg_man_output[180] = readOnlyReg(0);
    rg_man_output[181] = readOnlyReg(2);
    rg_man_output[182] = readOnlyReg(0);
    rg_man_output[183] = readOnlyReg(0);
    rg_man_output[184] = readOnlyReg(2);
    rg_man_output[185] = readOnlyReg(0);
    rg_man_output[186] = readOnlyReg(0);
    rg_man_output[187] = readOnlyReg(2);
    rg_man_output[188] = readOnlyReg(0);
    rg_man_output[189] = readOnlyReg(0);
    rg_man_output[190] = readOnlyReg(2);
    rg_man_output[191] = readOnlyReg(0);
    rg_man_output[192] = readOnlyReg(0);
    rg_man_output[193] = readOnlyReg(2);
    rg_man_output[194] = readOnlyReg(0);
    rg_man_output[195] = readOnlyReg(0);
    rg_man_output[196] = readOnlyReg(2);
    rg_man_output[197] = readOnlyReg(0);
    rg_man_output[198] = readOnlyReg(0);
    rg_man_output[199] = readOnlyReg(2);
    rg_man_output[200] = readOnlyReg(0);
    rg_man_output[201] = readOnlyReg(0);
    rg_man_output[202] = readOnlyReg(2);
    rg_man_output[203] = readOnlyReg(0);
    rg_man_output[204] = readOnlyReg(0);
    rg_man_output[205] = readOnlyReg(2);
    rg_man_output[206] = readOnlyReg(0);
    rg_man_output[207] = readOnlyReg(0);
    rg_man_output[208] = readOnlyReg(2);
    rg_man_output[209] = readOnlyReg(0);
    rg_man_output[210] = readOnlyReg(0);
    rg_man_output[211] = readOnlyReg(2);
    rg_man_output[212] = readOnlyReg(0);
    rg_man_output[213] = readOnlyReg(0);
    rg_man_output[214] = readOnlyReg(2);
    rg_man_output[215] = readOnlyReg(0);
    rg_man_output[216] = readOnlyReg(0);
    rg_man_output[217] = readOnlyReg(2);
    rg_man_output[218] = readOnlyReg(0);
    rg_man_output[219] = readOnlyReg(0);
    rg_man_output[220] = readOnlyReg(2);
    rg_man_output[221] = readOnlyReg(0);
    rg_man_output[222] = readOnlyReg(0);
    rg_man_output[223] = readOnlyReg(2);
    rg_man_output[224] = readOnlyReg(0);
    rg_man_output[225] = readOnlyReg(0);
    rg_man_output[226] = readOnlyReg(2);
    rg_man_output[227] = readOnlyReg(0);
    rg_man_output[228] = readOnlyReg(0);
    rg_man_output[229] = readOnlyReg(2);
    rg_man_output[230] = readOnlyReg(0);
    rg_man_output[231] = readOnlyReg(0);
    rg_man_output[232] = readOnlyReg(2);
    rg_man_output[233] = readOnlyReg(0);
    rg_man_output[234] = readOnlyReg(0);
    rg_man_output[235] = readOnlyReg(2);
    rg_man_output[236] = readOnlyReg(0);
    rg_man_output[237] = readOnlyReg(0);
    rg_man_output[238] = readOnlyReg(2);
    rg_man_output[239] = readOnlyReg(0);
    rg_man_output[240] = readOnlyReg(0);
    rg_man_output[241] = readOnlyReg(2);
    rg_man_output[242] = readOnlyReg(0);
    rg_man_output[243] = readOnlyReg(0);
    rg_man_output[244] = readOnlyReg(2);
    rg_man_output[245] = readOnlyReg(0);
    rg_man_output[246] = readOnlyReg(0);
    rg_man_output[247] = readOnlyReg(2);
    rg_man_output[248] = readOnlyReg(0);
    rg_man_output[249] = readOnlyReg(0);
    rg_man_output[250] = readOnlyReg(2);
    rg_man_output[251] = readOnlyReg(0);
    rg_man_output[252] = readOnlyReg(0);
    rg_man_output[253] = readOnlyReg(2);
    rg_man_output[254] = readOnlyReg(0);
    rg_man_output[255] = readOnlyReg(0);
    rg_man_output[256] = readOnlyReg(2);
    rg_man_output[257] = readOnlyReg(0);
    rg_man_output[258] = readOnlyReg(0);
    rg_man_output[259] = readOnlyReg(2);
    rg_man_output[260] = readOnlyReg(0);
    rg_man_output[261] = readOnlyReg(0);
    rg_man_output[262] = readOnlyReg(2);
    rg_man_output[263] = readOnlyReg(0);
    rg_man_output[264] = readOnlyReg(0);
    rg_man_output[265] = readOnlyReg(2);
    rg_man_output[266] = readOnlyReg(0);
    rg_man_output[267] = readOnlyReg(0);
    rg_man_output[268] = readOnlyReg(2);
    rg_man_output[269] = readOnlyReg(0);
    rg_man_output[270] = readOnlyReg(0);
    rg_man_output[271] = readOnlyReg(2);
    rg_man_output[272] = readOnlyReg(0);
    rg_man_output[273] = readOnlyReg(0);
    rg_man_output[274] = readOnlyReg(2);
    rg_man_output[275] = readOnlyReg(0);
    rg_man_output[276] = readOnlyReg(0);
    rg_man_output[277] = readOnlyReg(2);
    rg_man_output[278] = readOnlyReg(0);
    rg_man_output[279] = readOnlyReg(0);
    rg_man_output[280] = readOnlyReg(2);
    rg_man_output[281] = readOnlyReg(0);
    rg_man_output[282] = readOnlyReg(0);
    rg_man_output[283] = readOnlyReg(2);
    rg_man_output[284] = readOnlyReg(0);
    rg_man_output[285] = readOnlyReg(0);
    rg_man_output[286] = readOnlyReg(2);
    rg_man_output[287] = readOnlyReg(0);
    rg_man_output[288] = readOnlyReg(0);
    rg_man_output[289] = readOnlyReg(2);
    rg_man_output[290] = readOnlyReg(0);
    rg_man_output[291] = readOnlyReg(0);
    rg_man_output[292] = readOnlyReg(2);
    rg_man_output[293] = readOnlyReg(0);
    rg_man_output[294] = readOnlyReg(0);
    rg_man_output[295] = readOnlyReg(2);
    rg_man_output[296] = readOnlyReg(0);
    rg_man_output[297] = readOnlyReg(0);
    rg_man_output[298] = readOnlyReg(2);
    rg_man_output[299] = readOnlyReg(0);
    rg_man_output[300] = readOnlyReg(0);
    rg_man_output[301] = readOnlyReg(2);
    rg_man_output[302] = readOnlyReg(0);
    rg_man_output[303] = readOnlyReg(0);
    rg_man_output[304] = readOnlyReg(2);
    rg_man_output[305] = readOnlyReg(0);
    rg_man_output[306] = readOnlyReg(0);
    rg_man_output[307] = readOnlyReg(2);
    rg_man_output[308] = readOnlyReg(0);
    rg_man_output[309] = readOnlyReg(0);
    rg_man_output[310] = readOnlyReg(2);
    rg_man_output[311] = readOnlyReg(0);
    rg_man_output[312] = readOnlyReg(0);
    rg_man_output[313] = readOnlyReg(2);
    rg_man_output[314] = readOnlyReg(0);
    rg_man_output[315] = readOnlyReg(0);
    rg_man_output[316] = readOnlyReg(2);
    rg_man_output[317] = readOnlyReg(0);
    rg_man_output[318] = readOnlyReg(0);
    rg_man_output[319] = readOnlyReg(2);
    rg_man_output[320] = readOnlyReg(0);
    rg_man_output[321] = readOnlyReg(0);
    rg_man_output[322] = readOnlyReg(2);
    rg_man_output[323] = readOnlyReg(0);
    rg_man_output[324] = readOnlyReg(0);
    rg_man_output[325] = readOnlyReg(2);
    rg_man_output[326] = readOnlyReg(0);
    rg_man_output[327] = readOnlyReg(0);
    rg_man_output[328] = readOnlyReg(2);
    rg_man_output[329] = readOnlyReg(0);
    rg_man_output[330] = readOnlyReg(0);
    rg_man_output[331] = readOnlyReg(2);
    rg_man_output[332] = readOnlyReg(0);
    rg_man_output[333] = readOnlyReg(0);
    rg_man_output[334] = readOnlyReg(2);
    rg_man_output[335] = readOnlyReg(0);
    rg_man_output[336] = readOnlyReg(0);
    rg_man_output[337] = readOnlyReg(2);
    rg_man_output[338] = readOnlyReg(0);
    rg_man_output[339] = readOnlyReg(0);
    rg_man_output[340] = readOnlyReg(2);
    rg_man_output[341] = readOnlyReg(0);
    rg_man_output[342] = readOnlyReg(0);
    rg_man_output[343] = readOnlyReg(2);
    rg_man_output[344] = readOnlyReg(0);
    rg_man_output[345] = readOnlyReg(0);
    rg_man_output[346] = readOnlyReg(2);
    rg_man_output[347] = readOnlyReg(0);
    rg_man_output[348] = readOnlyReg(0);
    rg_man_output[349] = readOnlyReg(2);

    Reg#(Int#(7)) rg_exp_output[350];
    rg_exp_output[0] = readOnlyReg(-53);
    rg_exp_output[1] = readOnlyReg(-53);
    rg_exp_output[2] = readOnlyReg(-53);
    rg_exp_output[3] = readOnlyReg(-52);
    rg_exp_output[4] = readOnlyReg(-51);
    rg_exp_output[5] = readOnlyReg(-52);
    rg_exp_output[6] = readOnlyReg(-51);
    rg_exp_output[7] = readOnlyReg(-50);
    rg_exp_output[8] = readOnlyReg(-51);
    rg_exp_output[9] = readOnlyReg(-50);
    rg_exp_output[10] = readOnlyReg(-49);
    rg_exp_output[11] = readOnlyReg(-50);
    rg_exp_output[12] = readOnlyReg(-49);
    rg_exp_output[13] = readOnlyReg(-48);
    rg_exp_output[14] = readOnlyReg(-49);
    rg_exp_output[15] = readOnlyReg(-48);
    rg_exp_output[16] = readOnlyReg(-47);
    rg_exp_output[17] = readOnlyReg(-48);
    rg_exp_output[18] = readOnlyReg(-47);
    rg_exp_output[19] = readOnlyReg(-46);
    rg_exp_output[20] = readOnlyReg(-47);
    rg_exp_output[21] = readOnlyReg(-46);
    rg_exp_output[22] = readOnlyReg(-45);
    rg_exp_output[23] = readOnlyReg(-46);
    rg_exp_output[24] = readOnlyReg(-45);
    rg_exp_output[25] = readOnlyReg(-44);
    rg_exp_output[26] = readOnlyReg(-45);
    rg_exp_output[27] = readOnlyReg(-44);
    rg_exp_output[28] = readOnlyReg(-43);
    rg_exp_output[29] = readOnlyReg(-44);
    rg_exp_output[30] = readOnlyReg(-43);
    rg_exp_output[31] = readOnlyReg(-42);
    rg_exp_output[32] = readOnlyReg(-43);
    rg_exp_output[33] = readOnlyReg(-42);
    rg_exp_output[34] = readOnlyReg(-41);
    rg_exp_output[35] = readOnlyReg(-42);
    rg_exp_output[36] = readOnlyReg(-41);
    rg_exp_output[37] = readOnlyReg(-40);
    rg_exp_output[38] = readOnlyReg(-41);
    rg_exp_output[39] = readOnlyReg(-40);
    rg_exp_output[40] = readOnlyReg(-39);
    rg_exp_output[41] = readOnlyReg(-40);
    rg_exp_output[42] = readOnlyReg(-39);
    rg_exp_output[43] = readOnlyReg(-38);
    rg_exp_output[44] = readOnlyReg(-39);
    rg_exp_output[45] = readOnlyReg(-38);
    rg_exp_output[46] = readOnlyReg(-37);
    rg_exp_output[47] = readOnlyReg(-38);
    rg_exp_output[48] = readOnlyReg(-37);
    rg_exp_output[49] = readOnlyReg(-36);
    rg_exp_output[50] = readOnlyReg(-37);
    rg_exp_output[51] = readOnlyReg(-36);
    rg_exp_output[52] = readOnlyReg(-35);
    rg_exp_output[53] = readOnlyReg(-36);
    rg_exp_output[54] = readOnlyReg(-35);
    rg_exp_output[55] = readOnlyReg(-34);
    rg_exp_output[56] = readOnlyReg(-35);
    rg_exp_output[57] = readOnlyReg(-34);
    rg_exp_output[58] = readOnlyReg(-33);
    rg_exp_output[59] = readOnlyReg(-34);
    rg_exp_output[60] = readOnlyReg(-33);
    rg_exp_output[61] = readOnlyReg(-32);
    rg_exp_output[62] = readOnlyReg(-33);
    rg_exp_output[63] = readOnlyReg(-32);
    rg_exp_output[64] = readOnlyReg(-31);
    rg_exp_output[65] = readOnlyReg(-32);
    rg_exp_output[66] = readOnlyReg(-31);
    rg_exp_output[67] = readOnlyReg(-30);
    rg_exp_output[68] = readOnlyReg(-31);
    rg_exp_output[69] = readOnlyReg(-30);
    rg_exp_output[70] = readOnlyReg(-29);
    rg_exp_output[71] = readOnlyReg(-30);
    rg_exp_output[72] = readOnlyReg(-29);
    rg_exp_output[73] = readOnlyReg(-28);
    rg_exp_output[74] = readOnlyReg(-29);
    rg_exp_output[75] = readOnlyReg(-28);
    rg_exp_output[76] = readOnlyReg(-27);
    rg_exp_output[77] = readOnlyReg(-28);
    rg_exp_output[78] = readOnlyReg(-27);
    rg_exp_output[79] = readOnlyReg(-26);
    rg_exp_output[80] = readOnlyReg(-27);
    rg_exp_output[81] = readOnlyReg(-26);
    rg_exp_output[82] = readOnlyReg(-25);
    rg_exp_output[83] = readOnlyReg(-26);
    rg_exp_output[84] = readOnlyReg(-25);
    rg_exp_output[85] = readOnlyReg(-24);
    rg_exp_output[86] = readOnlyReg(-25);
    rg_exp_output[87] = readOnlyReg(-24);
    rg_exp_output[88] = readOnlyReg(-23);
    rg_exp_output[89] = readOnlyReg(-24);
    rg_exp_output[90] = readOnlyReg(-23);
    rg_exp_output[91] = readOnlyReg(-22);
    rg_exp_output[92] = readOnlyReg(-23);
    rg_exp_output[93] = readOnlyReg(-22);
    rg_exp_output[94] = readOnlyReg(-21);
    rg_exp_output[95] = readOnlyReg(-22);
    rg_exp_output[96] = readOnlyReg(-21);
    rg_exp_output[97] = readOnlyReg(-20);
    rg_exp_output[98] = readOnlyReg(-21);
    rg_exp_output[99] = readOnlyReg(-20);
    rg_exp_output[100] = readOnlyReg(-19);
    rg_exp_output[101] = readOnlyReg(-20);
    rg_exp_output[102] = readOnlyReg(-19);
    rg_exp_output[103] = readOnlyReg(-18);
    rg_exp_output[104] = readOnlyReg(-19);
    rg_exp_output[105] = readOnlyReg(-18);
    rg_exp_output[106] = readOnlyReg(-17);
    rg_exp_output[107] = readOnlyReg(-18);
    rg_exp_output[108] = readOnlyReg(-17);
    rg_exp_output[109] = readOnlyReg(-16);
    rg_exp_output[110] = readOnlyReg(-17);
    rg_exp_output[111] = readOnlyReg(-16);
    rg_exp_output[112] = readOnlyReg(-15);
    rg_exp_output[113] = readOnlyReg(-16);
    rg_exp_output[114] = readOnlyReg(-15);
    rg_exp_output[115] = readOnlyReg(-14);
    rg_exp_output[116] = readOnlyReg(-15);
    rg_exp_output[117] = readOnlyReg(-14);
    rg_exp_output[118] = readOnlyReg(-13);
    rg_exp_output[119] = readOnlyReg(-14);
    rg_exp_output[120] = readOnlyReg(-13);
    rg_exp_output[121] = readOnlyReg(-12);
    rg_exp_output[122] = readOnlyReg(-13);
    rg_exp_output[123] = readOnlyReg(-12);
    rg_exp_output[124] = readOnlyReg(-11);
    rg_exp_output[125] = readOnlyReg(-12);
    rg_exp_output[126] = readOnlyReg(-11);
    rg_exp_output[127] = readOnlyReg(-10);
    rg_exp_output[128] = readOnlyReg(-11);
    rg_exp_output[129] = readOnlyReg(-10);
    rg_exp_output[130] = readOnlyReg(-9);
    rg_exp_output[131] = readOnlyReg(-10);
    rg_exp_output[132] = readOnlyReg(-9);
    rg_exp_output[133] = readOnlyReg(-8);
    rg_exp_output[134] = readOnlyReg(-9);
    rg_exp_output[135] = readOnlyReg(-8);
    rg_exp_output[136] = readOnlyReg(-7);
    rg_exp_output[137] = readOnlyReg(-8);
    rg_exp_output[138] = readOnlyReg(-7);
    rg_exp_output[139] = readOnlyReg(-6);
    rg_exp_output[140] = readOnlyReg(-7);
    rg_exp_output[141] = readOnlyReg(-6);
    rg_exp_output[142] = readOnlyReg(-5);
    rg_exp_output[143] = readOnlyReg(-6);
    rg_exp_output[144] = readOnlyReg(-5);
    rg_exp_output[145] = readOnlyReg(-4);
    rg_exp_output[146] = readOnlyReg(-5);
    rg_exp_output[147] = readOnlyReg(-4);
    rg_exp_output[148] = readOnlyReg(-3);
    rg_exp_output[149] = readOnlyReg(-4);
    rg_exp_output[150] = readOnlyReg(-3);
    rg_exp_output[151] = readOnlyReg(-2);
    rg_exp_output[152] = readOnlyReg(-3);
    rg_exp_output[153] = readOnlyReg(-2);
    rg_exp_output[154] = readOnlyReg(-1);
    rg_exp_output[155] = readOnlyReg(-2);
    rg_exp_output[156] = readOnlyReg(-1);
    rg_exp_output[157] = readOnlyReg(-1);
    rg_exp_output[158] = readOnlyReg(0);
    rg_exp_output[159] = readOnlyReg(0);
    rg_exp_output[160] = readOnlyReg(0);
    rg_exp_output[161] = readOnlyReg(0);
    rg_exp_output[162] = readOnlyReg(0);
    rg_exp_output[163] = readOnlyReg(0);
    rg_exp_output[164] = readOnlyReg(0);
    rg_exp_output[165] = readOnlyReg(-62);
    rg_exp_output[166] = readOnlyReg(-62);
    rg_exp_output[167] = readOnlyReg(-62);
    rg_exp_output[168] = readOnlyReg(-61);
    rg_exp_output[169] = readOnlyReg(-61);
    rg_exp_output[170] = readOnlyReg(-61);
    rg_exp_output[171] = readOnlyReg(-60);
    rg_exp_output[172] = readOnlyReg(-60);
    rg_exp_output[173] = readOnlyReg(-60);
    rg_exp_output[174] = readOnlyReg(-59);
    rg_exp_output[175] = readOnlyReg(-59);
    rg_exp_output[176] = readOnlyReg(-59);
    rg_exp_output[177] = readOnlyReg(-58);
    rg_exp_output[178] = readOnlyReg(-58);
    rg_exp_output[179] = readOnlyReg(-58);
    rg_exp_output[180] = readOnlyReg(-57);
    rg_exp_output[181] = readOnlyReg(-57);
    rg_exp_output[182] = readOnlyReg(-57);
    rg_exp_output[183] = readOnlyReg(-56);
    rg_exp_output[184] = readOnlyReg(-56);
    rg_exp_output[185] = readOnlyReg(-56);
    rg_exp_output[186] = readOnlyReg(-55);
    rg_exp_output[187] = readOnlyReg(-55);
    rg_exp_output[188] = readOnlyReg(-55);
    rg_exp_output[189] = readOnlyReg(-54);
    rg_exp_output[190] = readOnlyReg(-54);
    rg_exp_output[191] = readOnlyReg(-54);
    rg_exp_output[192] = readOnlyReg(-53);
    rg_exp_output[193] = readOnlyReg(-53);
    rg_exp_output[194] = readOnlyReg(-53);
    rg_exp_output[195] = readOnlyReg(-52);
    rg_exp_output[196] = readOnlyReg(-52);
    rg_exp_output[197] = readOnlyReg(-52);
    rg_exp_output[198] = readOnlyReg(-51);
    rg_exp_output[199] = readOnlyReg(-51);
    rg_exp_output[200] = readOnlyReg(-51);
    rg_exp_output[201] = readOnlyReg(-50);
    rg_exp_output[202] = readOnlyReg(-50);
    rg_exp_output[203] = readOnlyReg(-50);
    rg_exp_output[204] = readOnlyReg(-49);
    rg_exp_output[205] = readOnlyReg(-49);
    rg_exp_output[206] = readOnlyReg(-49);
    rg_exp_output[207] = readOnlyReg(-48);
    rg_exp_output[208] = readOnlyReg(-48);
    rg_exp_output[209] = readOnlyReg(-48);
    rg_exp_output[210] = readOnlyReg(-47);
    rg_exp_output[211] = readOnlyReg(-47);
    rg_exp_output[212] = readOnlyReg(-47);
    rg_exp_output[213] = readOnlyReg(-46);
    rg_exp_output[214] = readOnlyReg(-46);
    rg_exp_output[215] = readOnlyReg(-46);
    rg_exp_output[216] = readOnlyReg(-45);
    rg_exp_output[217] = readOnlyReg(-45);
    rg_exp_output[218] = readOnlyReg(-45);
    rg_exp_output[219] = readOnlyReg(-44);
    rg_exp_output[220] = readOnlyReg(-44);
    rg_exp_output[221] = readOnlyReg(-44);
    rg_exp_output[222] = readOnlyReg(-43);
    rg_exp_output[223] = readOnlyReg(-43);
    rg_exp_output[224] = readOnlyReg(-43);
    rg_exp_output[225] = readOnlyReg(-42);
    rg_exp_output[226] = readOnlyReg(-42);
    rg_exp_output[227] = readOnlyReg(-42);
    rg_exp_output[228] = readOnlyReg(-41);
    rg_exp_output[229] = readOnlyReg(-41);
    rg_exp_output[230] = readOnlyReg(-41);
    rg_exp_output[231] = readOnlyReg(-40);
    rg_exp_output[232] = readOnlyReg(-40);
    rg_exp_output[233] = readOnlyReg(-40);
    rg_exp_output[234] = readOnlyReg(-39);
    rg_exp_output[235] = readOnlyReg(-39);
    rg_exp_output[236] = readOnlyReg(-39);
    rg_exp_output[237] = readOnlyReg(-38);
    rg_exp_output[238] = readOnlyReg(-38);
    rg_exp_output[239] = readOnlyReg(-38);
    rg_exp_output[240] = readOnlyReg(-37);
    rg_exp_output[241] = readOnlyReg(-37);
    rg_exp_output[242] = readOnlyReg(-37);
    rg_exp_output[243] = readOnlyReg(-36);
    rg_exp_output[244] = readOnlyReg(-36);
    rg_exp_output[245] = readOnlyReg(-36);
    rg_exp_output[246] = readOnlyReg(-35);
    rg_exp_output[247] = readOnlyReg(-35);
    rg_exp_output[248] = readOnlyReg(-35);
    rg_exp_output[249] = readOnlyReg(-34);
    rg_exp_output[250] = readOnlyReg(-34);
    rg_exp_output[251] = readOnlyReg(-34);
    rg_exp_output[252] = readOnlyReg(-33);
    rg_exp_output[253] = readOnlyReg(-33);
    rg_exp_output[254] = readOnlyReg(-33);
    rg_exp_output[255] = readOnlyReg(-32);
    rg_exp_output[256] = readOnlyReg(-32);
    rg_exp_output[257] = readOnlyReg(-32);
    rg_exp_output[258] = readOnlyReg(-31);
    rg_exp_output[259] = readOnlyReg(-31);
    rg_exp_output[260] = readOnlyReg(-31);
    rg_exp_output[261] = readOnlyReg(-30);
    rg_exp_output[262] = readOnlyReg(-30);
    rg_exp_output[263] = readOnlyReg(-30);
    rg_exp_output[264] = readOnlyReg(-29);
    rg_exp_output[265] = readOnlyReg(-29);
    rg_exp_output[266] = readOnlyReg(-29);
    rg_exp_output[267] = readOnlyReg(-28);
    rg_exp_output[268] = readOnlyReg(-28);
    rg_exp_output[269] = readOnlyReg(-28);
    rg_exp_output[270] = readOnlyReg(-27);
    rg_exp_output[271] = readOnlyReg(-27);
    rg_exp_output[272] = readOnlyReg(-27);
    rg_exp_output[273] = readOnlyReg(-26);
    rg_exp_output[274] = readOnlyReg(-26);
    rg_exp_output[275] = readOnlyReg(-26);
    rg_exp_output[276] = readOnlyReg(-25);
    rg_exp_output[277] = readOnlyReg(-25);
    rg_exp_output[278] = readOnlyReg(-25);
    rg_exp_output[279] = readOnlyReg(-24);
    rg_exp_output[280] = readOnlyReg(-24);
    rg_exp_output[281] = readOnlyReg(-24);
    rg_exp_output[282] = readOnlyReg(-23);
    rg_exp_output[283] = readOnlyReg(-23);
    rg_exp_output[284] = readOnlyReg(-23);
    rg_exp_output[285] = readOnlyReg(-22);
    rg_exp_output[286] = readOnlyReg(-22);
    rg_exp_output[287] = readOnlyReg(-22);
    rg_exp_output[288] = readOnlyReg(-21);
    rg_exp_output[289] = readOnlyReg(-21);
    rg_exp_output[290] = readOnlyReg(-21);
    rg_exp_output[291] = readOnlyReg(-20);
    rg_exp_output[292] = readOnlyReg(-20);
    rg_exp_output[293] = readOnlyReg(-20);
    rg_exp_output[294] = readOnlyReg(-19);
    rg_exp_output[295] = readOnlyReg(-19);
    rg_exp_output[296] = readOnlyReg(-19);
    rg_exp_output[297] = readOnlyReg(-18);
    rg_exp_output[298] = readOnlyReg(-18);
    rg_exp_output[299] = readOnlyReg(-18);
    rg_exp_output[300] = readOnlyReg(-17);
    rg_exp_output[301] = readOnlyReg(-17);
    rg_exp_output[302] = readOnlyReg(-17);
    rg_exp_output[303] = readOnlyReg(-16);
    rg_exp_output[304] = readOnlyReg(-16);
    rg_exp_output[305] = readOnlyReg(-16);
    rg_exp_output[306] = readOnlyReg(-15);
    rg_exp_output[307] = readOnlyReg(-15);
    rg_exp_output[308] = readOnlyReg(-15);
    rg_exp_output[309] = readOnlyReg(-14);
    rg_exp_output[310] = readOnlyReg(-14);
    rg_exp_output[311] = readOnlyReg(-14);
    rg_exp_output[312] = readOnlyReg(-13);
    rg_exp_output[313] = readOnlyReg(-13);
    rg_exp_output[314] = readOnlyReg(-13);
    rg_exp_output[315] = readOnlyReg(-12);
    rg_exp_output[316] = readOnlyReg(-12);
    rg_exp_output[317] = readOnlyReg(-12);
    rg_exp_output[318] = readOnlyReg(-11);
    rg_exp_output[319] = readOnlyReg(-11);
    rg_exp_output[320] = readOnlyReg(-11);
    rg_exp_output[321] = readOnlyReg(-10);
    rg_exp_output[322] = readOnlyReg(-10);
    rg_exp_output[323] = readOnlyReg(-10);
    rg_exp_output[324] = readOnlyReg(-9);
    rg_exp_output[325] = readOnlyReg(-9);
    rg_exp_output[326] = readOnlyReg(-9);
    rg_exp_output[327] = readOnlyReg(-8);
    rg_exp_output[328] = readOnlyReg(-8);
    rg_exp_output[329] = readOnlyReg(-8);
    rg_exp_output[330] = readOnlyReg(-7);
    rg_exp_output[331] = readOnlyReg(-7);
    rg_exp_output[332] = readOnlyReg(-7);
    rg_exp_output[333] = readOnlyReg(-6);
    rg_exp_output[334] = readOnlyReg(-6);
    rg_exp_output[335] = readOnlyReg(-6);
    rg_exp_output[336] = readOnlyReg(-5);
    rg_exp_output[337] = readOnlyReg(-5);
    rg_exp_output[338] = readOnlyReg(-5);
    rg_exp_output[339] = readOnlyReg(-4);
    rg_exp_output[340] = readOnlyReg(-4);
    rg_exp_output[341] = readOnlyReg(-4);
    rg_exp_output[342] = readOnlyReg(-3);
    rg_exp_output[343] = readOnlyReg(-3);
    rg_exp_output[344] = readOnlyReg(-3);
    rg_exp_output[345] = readOnlyReg(-2);
    rg_exp_output[346] = readOnlyReg(-2);
    rg_exp_output[347] = readOnlyReg(-2);
    rg_exp_output[348] = readOnlyReg(-1);
    rg_exp_output[349] = readOnlyReg(-1);

    method Tuple2#(Int#(7), Bit#(2)) mv_sig_output(Bit#(2) exp, Bit#(2) man);
      Bit#(4) index = {exp, man};
      return tuple2(rg_exp_output[index], rg_man_output[index]);
    endmethod
  endmodule


endpackage
